magic
tech scmos
timestamp 1607438890
<< rotate >>
rect 2047 302 2058 304
rect 2233 302 2244 304
rect 156 167 167 169
rect 423 167 434 169
rect 690 167 701 169
rect 957 167 968 169
rect 1224 167 1235 169
rect 1491 167 1502 169
rect 1758 167 1769 169
rect 2044 167 2055 169
rect 133 163 135 165
rect 156 160 170 167
rect 400 163 402 165
rect 423 160 437 167
rect 667 163 669 165
rect 690 160 704 167
rect 934 163 936 165
rect 957 160 971 167
rect 1201 163 1203 165
rect 1224 160 1238 167
rect 1468 163 1470 165
rect 1491 160 1505 167
rect 1735 163 1737 165
rect 1758 160 1772 167
rect 2021 163 2023 165
rect 2044 160 2058 167
rect 159 158 170 160
rect 426 158 437 160
rect 693 158 704 160
rect 960 158 971 160
rect 1227 158 1238 160
rect 1494 158 1505 160
rect 1761 158 1772 160
rect 2047 158 2058 160
rect 156 23 167 25
rect 423 23 434 25
rect 690 23 701 25
rect 957 23 968 25
rect 1224 23 1235 25
rect 1491 23 1502 25
rect 1758 23 1769 25
rect 2044 23 2055 25
rect 133 19 135 21
rect 156 16 170 23
rect 400 19 402 21
rect 423 16 437 23
rect 667 19 669 21
rect 690 16 704 23
rect 934 19 936 21
rect 957 16 971 23
rect 1201 19 1203 21
rect 1224 16 1238 23
rect 1468 19 1470 21
rect 1491 16 1505 23
rect 1735 19 1737 21
rect 1758 16 1772 23
rect 2021 19 2023 21
rect 2044 16 2058 23
rect 159 14 170 16
rect 426 14 437 16
rect 693 14 704 16
rect 960 14 971 16
rect 1227 14 1238 16
rect 1494 14 1505 16
rect 1761 14 1772 16
rect 2047 14 2058 16
rect 156 -121 167 -119
rect 423 -121 434 -119
rect 690 -121 701 -119
rect 957 -121 968 -119
rect 1224 -121 1235 -119
rect 1491 -121 1502 -119
rect 1758 -121 1769 -119
rect 2044 -121 2055 -119
rect 133 -125 135 -123
rect 156 -128 170 -121
rect 400 -125 402 -123
rect 423 -128 437 -121
rect 667 -125 669 -123
rect 690 -128 704 -121
rect 934 -125 936 -123
rect 957 -128 971 -121
rect 1201 -125 1203 -123
rect 1224 -128 1238 -121
rect 1468 -125 1470 -123
rect 1491 -128 1505 -121
rect 1735 -125 1737 -123
rect 1758 -128 1772 -121
rect 2021 -125 2023 -123
rect 2044 -128 2058 -121
rect 159 -130 170 -128
rect 426 -130 437 -128
rect 693 -130 704 -128
rect 960 -130 971 -128
rect 1227 -130 1238 -128
rect 1494 -130 1505 -128
rect 1761 -130 1772 -128
rect 2047 -130 2058 -128
rect 156 -265 167 -263
rect 423 -265 434 -263
rect 690 -265 701 -263
rect 957 -265 968 -263
rect 1224 -265 1235 -263
rect 1491 -265 1502 -263
rect 1758 -265 1769 -263
rect 2044 -265 2055 -263
rect 133 -269 135 -267
rect 156 -272 170 -265
rect 400 -269 402 -267
rect 423 -272 437 -265
rect 667 -269 669 -267
rect 690 -272 704 -265
rect 934 -269 936 -267
rect 957 -272 971 -265
rect 1201 -269 1203 -267
rect 1224 -272 1238 -265
rect 1468 -269 1470 -267
rect 1491 -272 1505 -265
rect 1735 -269 1737 -267
rect 1758 -272 1772 -265
rect 2021 -269 2023 -267
rect 2044 -272 2058 -265
rect 159 -274 170 -272
rect 426 -274 437 -272
rect 693 -274 704 -272
rect 960 -274 971 -272
rect 1227 -274 1238 -272
rect 2047 -274 2058 -272
<< ab >>
rect 6 290 263 304
rect 6 286 88 290
rect 90 286 260 290
rect 262 286 263 290
rect 6 178 263 286
rect 6 174 88 178
rect 90 174 260 178
rect 262 174 263 178
rect 6 146 263 174
rect 6 142 88 146
rect 90 142 260 146
rect 262 142 263 146
rect 6 34 263 142
rect 6 30 88 34
rect 90 30 260 34
rect 262 30 263 34
rect 6 2 263 30
rect 6 -2 88 2
rect 90 -2 260 2
rect 262 -2 263 2
rect 6 -110 263 -2
rect 6 -114 88 -110
rect 90 -114 260 -110
rect 262 -114 263 -110
rect 6 -142 263 -114
rect 6 -146 88 -142
rect 90 -146 260 -142
rect 262 -146 263 -142
rect 6 -254 263 -146
rect 6 -258 88 -254
rect 90 -258 260 -254
rect 262 -258 263 -254
rect 6 -272 263 -258
rect 265 193 306 304
rect 311 290 530 304
rect 311 286 355 290
rect 357 286 527 290
rect 529 286 530 290
rect 265 190 307 193
rect 265 49 306 190
rect 311 178 530 286
rect 311 174 355 178
rect 357 174 527 178
rect 529 174 530 178
rect 311 146 530 174
rect 311 142 355 146
rect 357 142 527 146
rect 529 142 530 146
rect 265 46 307 49
rect 265 -95 306 46
rect 311 34 530 142
rect 311 30 355 34
rect 357 30 527 34
rect 529 30 530 34
rect 311 2 530 30
rect 311 -2 355 2
rect 357 -2 527 2
rect 529 -2 530 2
rect 265 -98 307 -95
rect 265 -239 306 -98
rect 311 -110 530 -2
rect 311 -114 355 -110
rect 357 -114 527 -110
rect 529 -114 530 -110
rect 311 -142 530 -114
rect 311 -146 355 -142
rect 357 -146 527 -142
rect 529 -146 530 -142
rect 265 -242 307 -239
rect 265 -272 306 -242
rect 311 -254 530 -146
rect 311 -258 355 -254
rect 357 -258 527 -254
rect 529 -258 530 -254
rect 311 -272 530 -258
rect 532 193 573 304
rect 578 290 797 304
rect 578 286 622 290
rect 624 286 794 290
rect 796 286 797 290
rect 532 190 574 193
rect 532 49 573 190
rect 578 178 797 286
rect 578 174 622 178
rect 624 174 794 178
rect 796 174 797 178
rect 578 146 797 174
rect 578 142 622 146
rect 624 142 794 146
rect 796 142 797 146
rect 532 46 574 49
rect 532 -95 573 46
rect 578 34 797 142
rect 578 30 622 34
rect 624 30 794 34
rect 796 30 797 34
rect 578 2 797 30
rect 578 -2 622 2
rect 624 -2 794 2
rect 796 -2 797 2
rect 532 -98 574 -95
rect 532 -239 573 -98
rect 578 -110 797 -2
rect 578 -114 622 -110
rect 624 -114 794 -110
rect 796 -114 797 -110
rect 578 -142 797 -114
rect 578 -146 622 -142
rect 624 -146 794 -142
rect 796 -146 797 -142
rect 532 -242 574 -239
rect 532 -272 573 -242
rect 578 -254 797 -146
rect 578 -258 622 -254
rect 624 -258 794 -254
rect 796 -258 797 -254
rect 578 -272 797 -258
rect 799 193 840 304
rect 845 290 1064 304
rect 845 286 889 290
rect 891 286 1061 290
rect 1063 286 1064 290
rect 799 190 841 193
rect 799 49 840 190
rect 845 178 1064 286
rect 845 174 889 178
rect 891 174 1061 178
rect 1063 174 1064 178
rect 845 146 1064 174
rect 845 142 889 146
rect 891 142 1061 146
rect 1063 142 1064 146
rect 799 46 841 49
rect 799 -95 840 46
rect 845 34 1064 142
rect 845 30 889 34
rect 891 30 1061 34
rect 1063 30 1064 34
rect 845 2 1064 30
rect 845 -2 889 2
rect 891 -2 1061 2
rect 1063 -2 1064 2
rect 799 -98 841 -95
rect 799 -239 840 -98
rect 845 -110 1064 -2
rect 845 -114 889 -110
rect 891 -114 1061 -110
rect 1063 -114 1064 -110
rect 845 -142 1064 -114
rect 845 -146 889 -142
rect 891 -146 1061 -142
rect 1063 -146 1064 -142
rect 799 -242 841 -239
rect 799 -272 840 -242
rect 845 -254 1064 -146
rect 845 -258 889 -254
rect 891 -258 1061 -254
rect 1063 -258 1064 -254
rect 845 -272 1064 -258
rect 1066 193 1107 304
rect 1112 290 1331 304
rect 1112 286 1156 290
rect 1158 286 1328 290
rect 1330 286 1331 290
rect 1066 190 1108 193
rect 1066 49 1107 190
rect 1112 178 1331 286
rect 1112 174 1156 178
rect 1158 174 1328 178
rect 1330 174 1331 178
rect 1112 146 1331 174
rect 1112 142 1156 146
rect 1158 142 1328 146
rect 1330 142 1331 146
rect 1066 46 1108 49
rect 1066 -95 1107 46
rect 1112 34 1331 142
rect 1112 30 1156 34
rect 1158 30 1328 34
rect 1330 30 1331 34
rect 1112 2 1331 30
rect 1112 -2 1156 2
rect 1158 -2 1328 2
rect 1330 -2 1331 2
rect 1066 -98 1108 -95
rect 1066 -239 1107 -98
rect 1112 -110 1331 -2
rect 1112 -114 1156 -110
rect 1158 -114 1328 -110
rect 1330 -114 1331 -110
rect 1112 -142 1331 -114
rect 1112 -146 1156 -142
rect 1158 -146 1328 -142
rect 1330 -146 1331 -142
rect 1066 -242 1108 -239
rect 1066 -272 1107 -242
rect 1112 -254 1331 -146
rect 1112 -258 1156 -254
rect 1158 -258 1328 -254
rect 1330 -258 1331 -254
rect 1112 -272 1331 -258
rect 1333 193 1374 304
rect 1379 290 1598 304
rect 1379 286 1423 290
rect 1425 286 1595 290
rect 1597 286 1598 290
rect 1333 190 1375 193
rect 1333 49 1374 190
rect 1379 178 1598 286
rect 1379 174 1423 178
rect 1425 174 1595 178
rect 1597 174 1598 178
rect 1379 146 1598 174
rect 1379 142 1423 146
rect 1425 142 1595 146
rect 1597 142 1598 146
rect 1333 46 1375 49
rect 1333 -95 1374 46
rect 1379 34 1598 142
rect 1379 30 1423 34
rect 1425 30 1595 34
rect 1597 30 1598 34
rect 1379 2 1598 30
rect 1379 -2 1423 2
rect 1425 -2 1595 2
rect 1597 -2 1598 2
rect 1333 -98 1375 -95
rect 1333 -239 1374 -98
rect 1379 -110 1598 -2
rect 1379 -114 1423 -110
rect 1425 -114 1595 -110
rect 1597 -114 1598 -110
rect 1379 -142 1598 -114
rect 1379 -146 1423 -142
rect 1425 -146 1595 -142
rect 1597 -146 1598 -142
rect 1333 -242 1375 -239
rect 1333 -272 1374 -242
rect 1379 -254 1598 -146
rect 1379 -258 1423 -254
rect 1425 -258 1595 -254
rect 1597 -258 1598 -254
rect 1379 -272 1598 -258
rect 1600 193 1641 304
rect 1646 290 1865 304
rect 1646 286 1690 290
rect 1692 286 1862 290
rect 1864 286 1865 290
rect 1600 190 1642 193
rect 1600 49 1641 190
rect 1646 178 1865 286
rect 1646 174 1690 178
rect 1692 174 1862 178
rect 1864 174 1865 178
rect 1646 146 1865 174
rect 1646 142 1690 146
rect 1692 142 1862 146
rect 1864 142 1865 146
rect 1600 46 1642 49
rect 1600 -95 1641 46
rect 1646 34 1865 142
rect 1646 30 1690 34
rect 1692 30 1862 34
rect 1864 30 1865 34
rect 1646 2 1865 30
rect 1646 -2 1690 2
rect 1692 -2 1862 2
rect 1864 -2 1865 2
rect 1600 -98 1642 -95
rect 1600 -239 1641 -98
rect 1646 -110 1865 -2
rect 1646 -114 1690 -110
rect 1692 -114 1862 -110
rect 1864 -114 1865 -110
rect 1646 -142 1865 -114
rect 1646 -146 1690 -142
rect 1692 -146 1862 -142
rect 1864 -146 1865 -142
rect 1600 -242 1642 -239
rect 1600 -272 1641 -242
rect 1646 -254 1865 -146
rect 1646 -258 1690 -254
rect 1692 -258 1862 -254
rect 1864 -258 1865 -254
rect 1646 -272 1865 -258
rect 1867 193 1908 304
rect 1910 290 2151 304
rect 1910 286 1976 290
rect 1978 286 2148 290
rect 2150 286 2151 290
rect 1867 190 1909 193
rect 1867 49 1908 190
rect 1910 178 2151 286
rect 1910 174 1976 178
rect 1978 174 2148 178
rect 2150 174 2151 178
rect 1910 146 2151 174
rect 1910 142 1976 146
rect 1978 142 2148 146
rect 2150 142 2151 146
rect 1867 46 1909 49
rect 1867 -95 1908 46
rect 1910 34 2151 142
rect 1910 30 1976 34
rect 1978 30 2148 34
rect 2150 30 2151 34
rect 1910 2 2151 30
rect 1910 -2 1976 2
rect 1978 -2 2148 2
rect 2150 -2 2151 2
rect 1867 -98 1909 -95
rect 1867 -239 1908 -98
rect 1910 -110 2151 -2
rect 1910 -114 1976 -110
rect 1978 -114 2148 -110
rect 2150 -114 2151 -110
rect 1910 -142 2151 -114
rect 1910 -146 1976 -142
rect 1978 -146 2148 -142
rect 2150 -146 2151 -142
rect 1867 -242 1909 -239
rect 1867 -272 1908 -242
rect 1910 -254 2151 -146
rect 1910 -258 1976 -254
rect 1978 -258 2148 -254
rect 2150 -258 2151 -254
rect 1910 -272 2151 -258
rect 2153 193 2194 304
rect 2153 190 2195 193
rect 2153 49 2194 190
rect 2153 46 2195 49
rect 2153 -95 2194 46
rect 2153 -98 2195 -95
rect 2153 -239 2194 -98
rect 2153 -242 2195 -239
rect 2153 -272 2194 -242
rect 2197 -272 2261 304
rect 2265 -272 2329 304
<< nwell >>
rect 1 264 2332 309
rect 1 120 2332 200
rect 1 -24 2332 56
rect 1 -168 2332 -88
rect 1 -277 2332 -232
<< pwell >>
rect 1 200 2332 264
rect 1 56 2332 120
rect 1 -88 2332 -24
rect 1 -232 2332 -168
<< poly >>
rect 15 291 17 296
rect 25 291 27 296
rect 95 298 97 302
rect 35 289 37 293
rect 55 291 57 296
rect 65 291 67 296
rect 15 275 17 278
rect 11 273 17 275
rect 11 271 13 273
rect 15 271 17 273
rect 11 269 17 271
rect 15 256 17 269
rect 25 267 27 278
rect 75 289 77 293
rect 55 275 57 278
rect 51 273 57 275
rect 51 271 53 273
rect 55 271 57 273
rect 35 267 37 271
rect 51 269 57 271
rect 21 265 27 267
rect 21 263 23 265
rect 25 263 27 265
rect 21 261 27 263
rect 31 265 37 267
rect 31 263 33 265
rect 35 263 37 265
rect 31 261 37 263
rect 22 256 24 261
rect 35 256 37 261
rect 55 256 57 269
rect 65 267 67 278
rect 118 295 120 300
rect 125 295 127 300
rect 143 298 145 302
rect 153 298 155 302
rect 163 298 165 302
rect 185 298 187 302
rect 195 298 197 302
rect 205 298 207 302
rect 108 286 110 291
rect 75 267 77 271
rect 61 265 67 267
rect 61 263 63 265
rect 65 263 67 265
rect 61 261 67 263
rect 71 265 77 267
rect 71 263 73 265
rect 75 263 77 265
rect 71 261 77 263
rect 62 256 64 261
rect 75 256 77 261
rect 95 260 97 273
rect 108 270 110 273
rect 223 295 225 300
rect 230 295 232 300
rect 253 298 255 302
rect 274 298 276 302
rect 281 298 283 302
rect 240 286 242 291
rect 362 298 364 302
rect 294 288 296 293
rect 322 291 324 296
rect 332 291 334 296
rect 274 274 276 277
rect 240 270 242 273
rect 101 268 110 270
rect 101 266 103 268
rect 105 266 107 268
rect 118 267 120 270
rect 125 267 127 270
rect 143 267 145 270
rect 153 267 155 270
rect 163 267 165 270
rect 185 267 187 270
rect 195 267 197 270
rect 205 267 207 270
rect 223 267 225 270
rect 230 267 232 270
rect 240 268 249 270
rect 101 264 107 266
rect 95 258 101 260
rect 95 256 97 258
rect 99 256 101 258
rect 15 240 17 245
rect 22 240 24 245
rect 35 243 37 247
rect 95 254 101 256
rect 95 251 97 254
rect 105 251 107 264
rect 115 265 121 267
rect 115 263 117 265
rect 119 263 121 265
rect 115 261 121 263
rect 125 265 147 267
rect 125 263 136 265
rect 138 263 143 265
rect 145 263 147 265
rect 125 261 147 263
rect 151 265 157 267
rect 151 263 153 265
rect 155 263 157 265
rect 151 261 157 263
rect 161 265 167 267
rect 161 263 163 265
rect 165 263 167 265
rect 161 261 167 263
rect 183 265 189 267
rect 183 263 185 265
rect 187 263 189 265
rect 183 261 189 263
rect 193 265 199 267
rect 193 263 195 265
rect 197 263 199 265
rect 193 261 199 263
rect 203 265 225 267
rect 203 263 205 265
rect 207 263 212 265
rect 214 263 225 265
rect 203 261 225 263
rect 229 265 235 267
rect 229 263 231 265
rect 233 263 235 265
rect 229 261 235 263
rect 115 258 117 261
rect 125 258 127 261
rect 145 258 147 261
rect 152 258 154 261
rect 55 240 57 245
rect 62 240 64 245
rect 75 243 77 247
rect 95 234 97 238
rect 105 236 107 241
rect 115 239 117 244
rect 125 239 127 244
rect 163 252 165 261
rect 185 252 187 261
rect 196 258 198 261
rect 203 258 205 261
rect 223 258 225 261
rect 233 258 235 261
rect 243 266 245 268
rect 247 266 249 268
rect 243 264 249 266
rect 243 251 245 264
rect 253 260 255 273
rect 270 272 276 274
rect 270 270 272 272
rect 274 270 276 272
rect 270 268 276 270
rect 249 258 255 260
rect 274 258 276 268
rect 281 267 283 277
rect 342 289 344 293
rect 322 275 324 278
rect 318 273 324 275
rect 318 271 320 273
rect 322 271 324 273
rect 294 267 296 270
rect 318 269 324 271
rect 280 265 286 267
rect 280 263 282 265
rect 284 263 286 265
rect 280 261 286 263
rect 290 265 296 267
rect 290 263 292 265
rect 294 263 296 265
rect 290 261 296 263
rect 284 258 286 261
rect 294 258 296 261
rect 249 256 251 258
rect 253 256 255 258
rect 249 254 255 256
rect 253 251 255 254
rect 223 239 225 244
rect 233 239 235 244
rect 145 234 147 238
rect 152 234 154 238
rect 163 234 165 238
rect 185 234 187 238
rect 196 234 198 238
rect 203 234 205 238
rect 243 236 245 241
rect 274 247 276 252
rect 284 247 286 252
rect 322 256 324 269
rect 332 267 334 278
rect 385 295 387 300
rect 392 295 394 300
rect 410 298 412 302
rect 420 298 422 302
rect 430 298 432 302
rect 452 298 454 302
rect 462 298 464 302
rect 472 298 474 302
rect 375 286 377 291
rect 342 267 344 271
rect 328 265 334 267
rect 328 263 330 265
rect 332 263 334 265
rect 328 261 334 263
rect 338 265 344 267
rect 338 263 340 265
rect 342 263 344 265
rect 338 261 344 263
rect 329 256 331 261
rect 342 256 344 261
rect 362 260 364 273
rect 375 270 377 273
rect 490 295 492 300
rect 497 295 499 300
rect 520 298 522 302
rect 541 298 543 302
rect 548 298 550 302
rect 507 286 509 291
rect 629 298 631 302
rect 561 288 563 293
rect 589 291 591 296
rect 599 291 601 296
rect 541 274 543 277
rect 507 270 509 273
rect 368 268 377 270
rect 368 266 370 268
rect 372 266 374 268
rect 385 267 387 270
rect 392 267 394 270
rect 410 267 412 270
rect 420 267 422 270
rect 430 267 432 270
rect 452 267 454 270
rect 462 267 464 270
rect 472 267 474 270
rect 490 267 492 270
rect 497 267 499 270
rect 507 268 516 270
rect 368 264 374 266
rect 362 258 368 260
rect 362 256 364 258
rect 366 256 368 258
rect 294 244 296 249
rect 362 254 368 256
rect 362 251 364 254
rect 372 251 374 264
rect 382 265 388 267
rect 382 263 384 265
rect 386 263 388 265
rect 382 261 388 263
rect 392 265 414 267
rect 392 263 403 265
rect 405 263 410 265
rect 412 263 414 265
rect 392 261 414 263
rect 418 265 424 267
rect 418 263 420 265
rect 422 263 424 265
rect 418 261 424 263
rect 428 265 434 267
rect 428 263 430 265
rect 432 263 434 265
rect 428 261 434 263
rect 450 265 456 267
rect 450 263 452 265
rect 454 263 456 265
rect 450 261 456 263
rect 460 265 466 267
rect 460 263 462 265
rect 464 263 466 265
rect 460 261 466 263
rect 470 265 492 267
rect 470 263 472 265
rect 474 263 479 265
rect 481 263 492 265
rect 470 261 492 263
rect 496 265 502 267
rect 496 263 498 265
rect 500 263 502 265
rect 496 261 502 263
rect 382 258 384 261
rect 392 258 394 261
rect 412 258 414 261
rect 419 258 421 261
rect 322 240 324 245
rect 329 240 331 245
rect 253 234 255 238
rect 342 243 344 247
rect 362 234 364 238
rect 372 236 374 241
rect 382 239 384 244
rect 392 239 394 244
rect 430 252 432 261
rect 452 252 454 261
rect 463 258 465 261
rect 470 258 472 261
rect 490 258 492 261
rect 500 258 502 261
rect 510 266 512 268
rect 514 266 516 268
rect 510 264 516 266
rect 510 251 512 264
rect 520 260 522 273
rect 537 272 543 274
rect 537 270 539 272
rect 541 270 543 272
rect 537 268 543 270
rect 516 258 522 260
rect 541 258 543 268
rect 548 267 550 277
rect 609 289 611 293
rect 589 275 591 278
rect 585 273 591 275
rect 585 271 587 273
rect 589 271 591 273
rect 561 267 563 270
rect 585 269 591 271
rect 547 265 553 267
rect 547 263 549 265
rect 551 263 553 265
rect 547 261 553 263
rect 557 265 563 267
rect 557 263 559 265
rect 561 263 563 265
rect 557 261 563 263
rect 551 258 553 261
rect 561 258 563 261
rect 516 256 518 258
rect 520 256 522 258
rect 516 254 522 256
rect 520 251 522 254
rect 490 239 492 244
rect 500 239 502 244
rect 412 234 414 238
rect 419 234 421 238
rect 430 234 432 238
rect 452 234 454 238
rect 463 234 465 238
rect 470 234 472 238
rect 510 236 512 241
rect 541 247 543 252
rect 551 247 553 252
rect 589 256 591 269
rect 599 267 601 278
rect 652 295 654 300
rect 659 295 661 300
rect 677 298 679 302
rect 687 298 689 302
rect 697 298 699 302
rect 719 298 721 302
rect 729 298 731 302
rect 739 298 741 302
rect 642 286 644 291
rect 609 267 611 271
rect 595 265 601 267
rect 595 263 597 265
rect 599 263 601 265
rect 595 261 601 263
rect 605 265 611 267
rect 605 263 607 265
rect 609 263 611 265
rect 605 261 611 263
rect 596 256 598 261
rect 609 256 611 261
rect 629 260 631 273
rect 642 270 644 273
rect 757 295 759 300
rect 764 295 766 300
rect 787 298 789 302
rect 808 298 810 302
rect 815 298 817 302
rect 774 286 776 291
rect 896 298 898 302
rect 828 288 830 293
rect 856 291 858 296
rect 866 291 868 296
rect 808 274 810 277
rect 774 270 776 273
rect 635 268 644 270
rect 635 266 637 268
rect 639 266 641 268
rect 652 267 654 270
rect 659 267 661 270
rect 677 267 679 270
rect 687 267 689 270
rect 697 267 699 270
rect 719 267 721 270
rect 729 267 731 270
rect 739 267 741 270
rect 757 267 759 270
rect 764 267 766 270
rect 774 268 783 270
rect 635 264 641 266
rect 629 258 635 260
rect 629 256 631 258
rect 633 256 635 258
rect 561 244 563 249
rect 629 254 635 256
rect 629 251 631 254
rect 639 251 641 264
rect 649 265 655 267
rect 649 263 651 265
rect 653 263 655 265
rect 649 261 655 263
rect 659 265 681 267
rect 659 263 670 265
rect 672 263 677 265
rect 679 263 681 265
rect 659 261 681 263
rect 685 265 691 267
rect 685 263 687 265
rect 689 263 691 265
rect 685 261 691 263
rect 695 265 701 267
rect 695 263 697 265
rect 699 263 701 265
rect 695 261 701 263
rect 717 265 723 267
rect 717 263 719 265
rect 721 263 723 265
rect 717 261 723 263
rect 727 265 733 267
rect 727 263 729 265
rect 731 263 733 265
rect 727 261 733 263
rect 737 265 759 267
rect 737 263 739 265
rect 741 263 746 265
rect 748 263 759 265
rect 737 261 759 263
rect 763 265 769 267
rect 763 263 765 265
rect 767 263 769 265
rect 763 261 769 263
rect 649 258 651 261
rect 659 258 661 261
rect 679 258 681 261
rect 686 258 688 261
rect 589 240 591 245
rect 596 240 598 245
rect 520 234 522 238
rect 609 243 611 247
rect 629 234 631 238
rect 639 236 641 241
rect 649 239 651 244
rect 659 239 661 244
rect 697 252 699 261
rect 719 252 721 261
rect 730 258 732 261
rect 737 258 739 261
rect 757 258 759 261
rect 767 258 769 261
rect 777 266 779 268
rect 781 266 783 268
rect 777 264 783 266
rect 777 251 779 264
rect 787 260 789 273
rect 804 272 810 274
rect 804 270 806 272
rect 808 270 810 272
rect 804 268 810 270
rect 783 258 789 260
rect 808 258 810 268
rect 815 267 817 277
rect 876 289 878 293
rect 856 275 858 278
rect 852 273 858 275
rect 852 271 854 273
rect 856 271 858 273
rect 828 267 830 270
rect 852 269 858 271
rect 814 265 820 267
rect 814 263 816 265
rect 818 263 820 265
rect 814 261 820 263
rect 824 265 830 267
rect 824 263 826 265
rect 828 263 830 265
rect 824 261 830 263
rect 818 258 820 261
rect 828 258 830 261
rect 783 256 785 258
rect 787 256 789 258
rect 783 254 789 256
rect 787 251 789 254
rect 757 239 759 244
rect 767 239 769 244
rect 679 234 681 238
rect 686 234 688 238
rect 697 234 699 238
rect 719 234 721 238
rect 730 234 732 238
rect 737 234 739 238
rect 777 236 779 241
rect 808 247 810 252
rect 818 247 820 252
rect 856 256 858 269
rect 866 267 868 278
rect 919 295 921 300
rect 926 295 928 300
rect 944 298 946 302
rect 954 298 956 302
rect 964 298 966 302
rect 986 298 988 302
rect 996 298 998 302
rect 1006 298 1008 302
rect 909 286 911 291
rect 876 267 878 271
rect 862 265 868 267
rect 862 263 864 265
rect 866 263 868 265
rect 862 261 868 263
rect 872 265 878 267
rect 872 263 874 265
rect 876 263 878 265
rect 872 261 878 263
rect 863 256 865 261
rect 876 256 878 261
rect 896 260 898 273
rect 909 270 911 273
rect 1024 295 1026 300
rect 1031 295 1033 300
rect 1054 298 1056 302
rect 1075 298 1077 302
rect 1082 298 1084 302
rect 1041 286 1043 291
rect 1163 298 1165 302
rect 1095 288 1097 293
rect 1123 291 1125 296
rect 1133 291 1135 296
rect 1075 274 1077 277
rect 1041 270 1043 273
rect 902 268 911 270
rect 902 266 904 268
rect 906 266 908 268
rect 919 267 921 270
rect 926 267 928 270
rect 944 267 946 270
rect 954 267 956 270
rect 964 267 966 270
rect 986 267 988 270
rect 996 267 998 270
rect 1006 267 1008 270
rect 1024 267 1026 270
rect 1031 267 1033 270
rect 1041 268 1050 270
rect 902 264 908 266
rect 896 258 902 260
rect 896 256 898 258
rect 900 256 902 258
rect 828 244 830 249
rect 896 254 902 256
rect 896 251 898 254
rect 906 251 908 264
rect 916 265 922 267
rect 916 263 918 265
rect 920 263 922 265
rect 916 261 922 263
rect 926 265 948 267
rect 926 263 937 265
rect 939 263 944 265
rect 946 263 948 265
rect 926 261 948 263
rect 952 265 958 267
rect 952 263 954 265
rect 956 263 958 265
rect 952 261 958 263
rect 962 265 968 267
rect 962 263 964 265
rect 966 263 968 265
rect 962 261 968 263
rect 984 265 990 267
rect 984 263 986 265
rect 988 263 990 265
rect 984 261 990 263
rect 994 265 1000 267
rect 994 263 996 265
rect 998 263 1000 265
rect 994 261 1000 263
rect 1004 265 1026 267
rect 1004 263 1006 265
rect 1008 263 1013 265
rect 1015 263 1026 265
rect 1004 261 1026 263
rect 1030 265 1036 267
rect 1030 263 1032 265
rect 1034 263 1036 265
rect 1030 261 1036 263
rect 916 258 918 261
rect 926 258 928 261
rect 946 258 948 261
rect 953 258 955 261
rect 856 240 858 245
rect 863 240 865 245
rect 787 234 789 238
rect 876 243 878 247
rect 896 234 898 238
rect 906 236 908 241
rect 916 239 918 244
rect 926 239 928 244
rect 964 252 966 261
rect 986 252 988 261
rect 997 258 999 261
rect 1004 258 1006 261
rect 1024 258 1026 261
rect 1034 258 1036 261
rect 1044 266 1046 268
rect 1048 266 1050 268
rect 1044 264 1050 266
rect 1044 251 1046 264
rect 1054 260 1056 273
rect 1071 272 1077 274
rect 1071 270 1073 272
rect 1075 270 1077 272
rect 1071 268 1077 270
rect 1050 258 1056 260
rect 1075 258 1077 268
rect 1082 267 1084 277
rect 1143 289 1145 293
rect 1123 275 1125 278
rect 1119 273 1125 275
rect 1119 271 1121 273
rect 1123 271 1125 273
rect 1095 267 1097 270
rect 1119 269 1125 271
rect 1081 265 1087 267
rect 1081 263 1083 265
rect 1085 263 1087 265
rect 1081 261 1087 263
rect 1091 265 1097 267
rect 1091 263 1093 265
rect 1095 263 1097 265
rect 1091 261 1097 263
rect 1085 258 1087 261
rect 1095 258 1097 261
rect 1050 256 1052 258
rect 1054 256 1056 258
rect 1050 254 1056 256
rect 1054 251 1056 254
rect 1024 239 1026 244
rect 1034 239 1036 244
rect 946 234 948 238
rect 953 234 955 238
rect 964 234 966 238
rect 986 234 988 238
rect 997 234 999 238
rect 1004 234 1006 238
rect 1044 236 1046 241
rect 1075 247 1077 252
rect 1085 247 1087 252
rect 1123 256 1125 269
rect 1133 267 1135 278
rect 1186 295 1188 300
rect 1193 295 1195 300
rect 1211 298 1213 302
rect 1221 298 1223 302
rect 1231 298 1233 302
rect 1253 298 1255 302
rect 1263 298 1265 302
rect 1273 298 1275 302
rect 1176 286 1178 291
rect 1143 267 1145 271
rect 1129 265 1135 267
rect 1129 263 1131 265
rect 1133 263 1135 265
rect 1129 261 1135 263
rect 1139 265 1145 267
rect 1139 263 1141 265
rect 1143 263 1145 265
rect 1139 261 1145 263
rect 1130 256 1132 261
rect 1143 256 1145 261
rect 1163 260 1165 273
rect 1176 270 1178 273
rect 1291 295 1293 300
rect 1298 295 1300 300
rect 1321 298 1323 302
rect 1342 298 1344 302
rect 1349 298 1351 302
rect 1308 286 1310 291
rect 1430 298 1432 302
rect 1362 288 1364 293
rect 1390 291 1392 296
rect 1400 291 1402 296
rect 1342 274 1344 277
rect 1308 270 1310 273
rect 1169 268 1178 270
rect 1169 266 1171 268
rect 1173 266 1175 268
rect 1186 267 1188 270
rect 1193 267 1195 270
rect 1211 267 1213 270
rect 1221 267 1223 270
rect 1231 267 1233 270
rect 1253 267 1255 270
rect 1263 267 1265 270
rect 1273 267 1275 270
rect 1291 267 1293 270
rect 1298 267 1300 270
rect 1308 268 1317 270
rect 1169 264 1175 266
rect 1163 258 1169 260
rect 1163 256 1165 258
rect 1167 256 1169 258
rect 1095 244 1097 249
rect 1163 254 1169 256
rect 1163 251 1165 254
rect 1173 251 1175 264
rect 1183 265 1189 267
rect 1183 263 1185 265
rect 1187 263 1189 265
rect 1183 261 1189 263
rect 1193 265 1215 267
rect 1193 263 1204 265
rect 1206 263 1211 265
rect 1213 263 1215 265
rect 1193 261 1215 263
rect 1219 265 1225 267
rect 1219 263 1221 265
rect 1223 263 1225 265
rect 1219 261 1225 263
rect 1229 265 1235 267
rect 1229 263 1231 265
rect 1233 263 1235 265
rect 1229 261 1235 263
rect 1251 265 1257 267
rect 1251 263 1253 265
rect 1255 263 1257 265
rect 1251 261 1257 263
rect 1261 265 1267 267
rect 1261 263 1263 265
rect 1265 263 1267 265
rect 1261 261 1267 263
rect 1271 265 1293 267
rect 1271 263 1273 265
rect 1275 263 1280 265
rect 1282 263 1293 265
rect 1271 261 1293 263
rect 1297 265 1303 267
rect 1297 263 1299 265
rect 1301 263 1303 265
rect 1297 261 1303 263
rect 1183 258 1185 261
rect 1193 258 1195 261
rect 1213 258 1215 261
rect 1220 258 1222 261
rect 1123 240 1125 245
rect 1130 240 1132 245
rect 1054 234 1056 238
rect 1143 243 1145 247
rect 1163 234 1165 238
rect 1173 236 1175 241
rect 1183 239 1185 244
rect 1193 239 1195 244
rect 1231 252 1233 261
rect 1253 252 1255 261
rect 1264 258 1266 261
rect 1271 258 1273 261
rect 1291 258 1293 261
rect 1301 258 1303 261
rect 1311 266 1313 268
rect 1315 266 1317 268
rect 1311 264 1317 266
rect 1311 251 1313 264
rect 1321 260 1323 273
rect 1338 272 1344 274
rect 1338 270 1340 272
rect 1342 270 1344 272
rect 1338 268 1344 270
rect 1317 258 1323 260
rect 1342 258 1344 268
rect 1349 267 1351 277
rect 1410 289 1412 293
rect 1390 275 1392 278
rect 1386 273 1392 275
rect 1386 271 1388 273
rect 1390 271 1392 273
rect 1362 267 1364 270
rect 1386 269 1392 271
rect 1348 265 1354 267
rect 1348 263 1350 265
rect 1352 263 1354 265
rect 1348 261 1354 263
rect 1358 265 1364 267
rect 1358 263 1360 265
rect 1362 263 1364 265
rect 1358 261 1364 263
rect 1352 258 1354 261
rect 1362 258 1364 261
rect 1317 256 1319 258
rect 1321 256 1323 258
rect 1317 254 1323 256
rect 1321 251 1323 254
rect 1291 239 1293 244
rect 1301 239 1303 244
rect 1213 234 1215 238
rect 1220 234 1222 238
rect 1231 234 1233 238
rect 1253 234 1255 238
rect 1264 234 1266 238
rect 1271 234 1273 238
rect 1311 236 1313 241
rect 1342 247 1344 252
rect 1352 247 1354 252
rect 1390 256 1392 269
rect 1400 267 1402 278
rect 1453 295 1455 300
rect 1460 295 1462 300
rect 1478 298 1480 302
rect 1488 298 1490 302
rect 1498 298 1500 302
rect 1520 298 1522 302
rect 1530 298 1532 302
rect 1540 298 1542 302
rect 1443 286 1445 291
rect 1410 267 1412 271
rect 1396 265 1402 267
rect 1396 263 1398 265
rect 1400 263 1402 265
rect 1396 261 1402 263
rect 1406 265 1412 267
rect 1406 263 1408 265
rect 1410 263 1412 265
rect 1406 261 1412 263
rect 1397 256 1399 261
rect 1410 256 1412 261
rect 1430 260 1432 273
rect 1443 270 1445 273
rect 1558 295 1560 300
rect 1565 295 1567 300
rect 1588 298 1590 302
rect 1609 298 1611 302
rect 1616 298 1618 302
rect 1575 286 1577 291
rect 1697 298 1699 302
rect 1629 288 1631 293
rect 1657 291 1659 296
rect 1667 291 1669 296
rect 1609 274 1611 277
rect 1575 270 1577 273
rect 1436 268 1445 270
rect 1436 266 1438 268
rect 1440 266 1442 268
rect 1453 267 1455 270
rect 1460 267 1462 270
rect 1478 267 1480 270
rect 1488 267 1490 270
rect 1498 267 1500 270
rect 1520 267 1522 270
rect 1530 267 1532 270
rect 1540 267 1542 270
rect 1558 267 1560 270
rect 1565 267 1567 270
rect 1575 268 1584 270
rect 1436 264 1442 266
rect 1430 258 1436 260
rect 1430 256 1432 258
rect 1434 256 1436 258
rect 1362 244 1364 249
rect 1430 254 1436 256
rect 1430 251 1432 254
rect 1440 251 1442 264
rect 1450 265 1456 267
rect 1450 263 1452 265
rect 1454 263 1456 265
rect 1450 261 1456 263
rect 1460 265 1482 267
rect 1460 263 1471 265
rect 1473 263 1478 265
rect 1480 263 1482 265
rect 1460 261 1482 263
rect 1486 265 1492 267
rect 1486 263 1488 265
rect 1490 263 1492 265
rect 1486 261 1492 263
rect 1496 265 1502 267
rect 1496 263 1498 265
rect 1500 263 1502 265
rect 1496 261 1502 263
rect 1518 265 1524 267
rect 1518 263 1520 265
rect 1522 263 1524 265
rect 1518 261 1524 263
rect 1528 265 1534 267
rect 1528 263 1530 265
rect 1532 263 1534 265
rect 1528 261 1534 263
rect 1538 265 1560 267
rect 1538 263 1540 265
rect 1542 263 1547 265
rect 1549 263 1560 265
rect 1538 261 1560 263
rect 1564 265 1570 267
rect 1564 263 1566 265
rect 1568 263 1570 265
rect 1564 261 1570 263
rect 1450 258 1452 261
rect 1460 258 1462 261
rect 1480 258 1482 261
rect 1487 258 1489 261
rect 1390 240 1392 245
rect 1397 240 1399 245
rect 1321 234 1323 238
rect 1410 243 1412 247
rect 1430 234 1432 238
rect 1440 236 1442 241
rect 1450 239 1452 244
rect 1460 239 1462 244
rect 1498 252 1500 261
rect 1520 252 1522 261
rect 1531 258 1533 261
rect 1538 258 1540 261
rect 1558 258 1560 261
rect 1568 258 1570 261
rect 1578 266 1580 268
rect 1582 266 1584 268
rect 1578 264 1584 266
rect 1578 251 1580 264
rect 1588 260 1590 273
rect 1605 272 1611 274
rect 1605 270 1607 272
rect 1609 270 1611 272
rect 1605 268 1611 270
rect 1584 258 1590 260
rect 1609 258 1611 268
rect 1616 267 1618 277
rect 1677 289 1679 293
rect 1657 275 1659 278
rect 1653 273 1659 275
rect 1653 271 1655 273
rect 1657 271 1659 273
rect 1629 267 1631 270
rect 1653 269 1659 271
rect 1615 265 1621 267
rect 1615 263 1617 265
rect 1619 263 1621 265
rect 1615 261 1621 263
rect 1625 265 1631 267
rect 1625 263 1627 265
rect 1629 263 1631 265
rect 1625 261 1631 263
rect 1619 258 1621 261
rect 1629 258 1631 261
rect 1584 256 1586 258
rect 1588 256 1590 258
rect 1584 254 1590 256
rect 1588 251 1590 254
rect 1558 239 1560 244
rect 1568 239 1570 244
rect 1480 234 1482 238
rect 1487 234 1489 238
rect 1498 234 1500 238
rect 1520 234 1522 238
rect 1531 234 1533 238
rect 1538 234 1540 238
rect 1578 236 1580 241
rect 1609 247 1611 252
rect 1619 247 1621 252
rect 1657 256 1659 269
rect 1667 267 1669 278
rect 1720 295 1722 300
rect 1727 295 1729 300
rect 1745 298 1747 302
rect 1755 298 1757 302
rect 1765 298 1767 302
rect 1787 298 1789 302
rect 1797 298 1799 302
rect 1807 298 1809 302
rect 1710 286 1712 291
rect 1677 267 1679 271
rect 1663 265 1669 267
rect 1663 263 1665 265
rect 1667 263 1669 265
rect 1663 261 1669 263
rect 1673 265 1679 267
rect 1673 263 1675 265
rect 1677 263 1679 265
rect 1673 261 1679 263
rect 1664 256 1666 261
rect 1677 256 1679 261
rect 1697 260 1699 273
rect 1710 270 1712 273
rect 1825 295 1827 300
rect 1832 295 1834 300
rect 1855 298 1857 302
rect 1876 298 1878 302
rect 1883 298 1885 302
rect 1842 286 1844 291
rect 1927 298 1929 302
rect 1896 288 1898 293
rect 1876 274 1878 277
rect 1842 270 1844 273
rect 1703 268 1712 270
rect 1703 266 1705 268
rect 1707 266 1709 268
rect 1720 267 1722 270
rect 1727 267 1729 270
rect 1745 267 1747 270
rect 1755 267 1757 270
rect 1765 267 1767 270
rect 1787 267 1789 270
rect 1797 267 1799 270
rect 1807 267 1809 270
rect 1825 267 1827 270
rect 1832 267 1834 270
rect 1842 268 1851 270
rect 1703 264 1709 266
rect 1697 258 1703 260
rect 1697 256 1699 258
rect 1701 256 1703 258
rect 1629 244 1631 249
rect 1697 254 1703 256
rect 1697 251 1699 254
rect 1707 251 1709 264
rect 1717 265 1723 267
rect 1717 263 1719 265
rect 1721 263 1723 265
rect 1717 261 1723 263
rect 1727 265 1749 267
rect 1727 263 1738 265
rect 1740 263 1745 265
rect 1747 263 1749 265
rect 1727 261 1749 263
rect 1753 265 1759 267
rect 1753 263 1755 265
rect 1757 263 1759 265
rect 1753 261 1759 263
rect 1763 265 1769 267
rect 1763 263 1765 265
rect 1767 263 1769 265
rect 1763 261 1769 263
rect 1785 265 1791 267
rect 1785 263 1787 265
rect 1789 263 1791 265
rect 1785 261 1791 263
rect 1795 265 1801 267
rect 1795 263 1797 265
rect 1799 263 1801 265
rect 1795 261 1801 263
rect 1805 265 1827 267
rect 1805 263 1807 265
rect 1809 263 1814 265
rect 1816 263 1827 265
rect 1805 261 1827 263
rect 1831 265 1837 267
rect 1831 263 1833 265
rect 1835 263 1837 265
rect 1831 261 1837 263
rect 1717 258 1719 261
rect 1727 258 1729 261
rect 1747 258 1749 261
rect 1754 258 1756 261
rect 1657 240 1659 245
rect 1664 240 1666 245
rect 1588 234 1590 238
rect 1677 243 1679 247
rect 1697 234 1699 238
rect 1707 236 1709 241
rect 1717 239 1719 244
rect 1727 239 1729 244
rect 1765 252 1767 261
rect 1787 252 1789 261
rect 1798 258 1800 261
rect 1805 258 1807 261
rect 1825 258 1827 261
rect 1835 258 1837 261
rect 1845 266 1847 268
rect 1849 266 1851 268
rect 1845 264 1851 266
rect 1845 251 1847 264
rect 1855 260 1857 273
rect 1872 272 1878 274
rect 1872 270 1874 272
rect 1876 270 1878 272
rect 1872 268 1878 270
rect 1851 258 1857 260
rect 1876 258 1878 268
rect 1883 267 1885 277
rect 1912 273 1918 275
rect 1912 271 1914 273
rect 1916 271 1918 273
rect 1963 298 1965 302
rect 1983 298 1985 302
rect 1943 289 1945 293
rect 1953 289 1955 293
rect 2006 295 2008 300
rect 2013 295 2015 300
rect 2031 298 2033 302
rect 2041 298 2043 302
rect 2051 298 2053 302
rect 2073 298 2075 302
rect 2083 298 2085 302
rect 2093 298 2095 302
rect 1996 286 1998 291
rect 1896 267 1898 270
rect 1912 269 1918 271
rect 1882 265 1888 267
rect 1882 263 1884 265
rect 1886 263 1888 265
rect 1882 261 1888 263
rect 1892 265 1898 267
rect 1916 268 1918 269
rect 1927 268 1929 271
rect 1943 268 1945 271
rect 1916 266 1929 268
rect 1935 266 1945 268
rect 1953 267 1955 271
rect 1963 268 1965 271
rect 1892 263 1894 265
rect 1896 263 1898 265
rect 1892 261 1898 263
rect 1886 258 1888 261
rect 1896 258 1898 261
rect 1919 258 1921 266
rect 1935 262 1937 266
rect 1928 260 1937 262
rect 1949 265 1955 267
rect 1949 263 1951 265
rect 1953 263 1955 265
rect 1949 261 1955 263
rect 1959 266 1965 268
rect 1959 264 1961 266
rect 1963 264 1965 266
rect 1959 262 1965 264
rect 1928 258 1930 260
rect 1932 258 1937 260
rect 1851 256 1853 258
rect 1855 256 1857 258
rect 1851 254 1857 256
rect 1855 251 1857 254
rect 1825 239 1827 244
rect 1835 239 1837 244
rect 1747 234 1749 238
rect 1754 234 1756 238
rect 1765 234 1767 238
rect 1787 234 1789 238
rect 1798 234 1800 238
rect 1805 234 1807 238
rect 1845 236 1847 241
rect 1876 247 1878 252
rect 1886 247 1888 252
rect 1928 256 1937 258
rect 1953 258 1955 261
rect 1935 253 1937 256
rect 1945 253 1947 257
rect 1953 256 1957 258
rect 1955 253 1957 256
rect 1962 253 1964 262
rect 1983 260 1985 273
rect 1996 270 1998 273
rect 2111 295 2113 300
rect 2118 295 2120 300
rect 2141 298 2143 302
rect 2162 298 2164 302
rect 2169 298 2171 302
rect 2128 286 2130 291
rect 2216 298 2218 302
rect 2223 298 2225 302
rect 2233 298 2235 302
rect 2240 298 2242 302
rect 2250 298 2252 302
rect 2284 298 2286 302
rect 2291 298 2293 302
rect 2301 298 2303 302
rect 2308 298 2310 302
rect 2318 298 2320 302
rect 2182 288 2184 293
rect 2162 274 2164 277
rect 2128 270 2130 273
rect 1989 268 1998 270
rect 1989 266 1991 268
rect 1993 266 1995 268
rect 2006 267 2008 270
rect 2013 267 2015 270
rect 2031 267 2033 270
rect 2041 267 2043 270
rect 2051 267 2053 270
rect 2073 267 2075 270
rect 2083 267 2085 270
rect 2093 267 2095 270
rect 2111 267 2113 270
rect 2118 267 2120 270
rect 2128 268 2137 270
rect 1989 264 1995 266
rect 1983 258 1989 260
rect 1983 256 1985 258
rect 1987 256 1989 258
rect 1983 254 1989 256
rect 1896 244 1898 249
rect 1919 246 1921 249
rect 1919 244 1924 246
rect 1855 234 1857 238
rect 1922 236 1924 244
rect 1935 240 1937 244
rect 1945 236 1947 244
rect 1983 251 1985 254
rect 1993 251 1995 264
rect 2003 265 2009 267
rect 2003 263 2005 265
rect 2007 263 2009 265
rect 2003 261 2009 263
rect 2013 265 2035 267
rect 2013 263 2024 265
rect 2026 263 2031 265
rect 2033 263 2035 265
rect 2013 261 2035 263
rect 2039 265 2045 267
rect 2039 263 2041 265
rect 2043 263 2045 265
rect 2039 261 2045 263
rect 2049 265 2055 267
rect 2049 263 2051 265
rect 2053 263 2055 265
rect 2049 261 2055 263
rect 2071 265 2077 267
rect 2071 263 2073 265
rect 2075 263 2077 265
rect 2071 261 2077 263
rect 2081 265 2087 267
rect 2081 263 2083 265
rect 2085 263 2087 265
rect 2081 261 2087 263
rect 2091 265 2113 267
rect 2091 263 2093 265
rect 2095 263 2100 265
rect 2102 263 2113 265
rect 2091 261 2113 263
rect 2117 265 2123 267
rect 2117 263 2119 265
rect 2121 263 2123 265
rect 2117 261 2123 263
rect 2003 258 2005 261
rect 2013 258 2015 261
rect 2033 258 2035 261
rect 2040 258 2042 261
rect 1955 236 1957 241
rect 1962 236 1964 241
rect 1922 234 1947 236
rect 1983 234 1985 238
rect 1993 236 1995 241
rect 2003 239 2005 244
rect 2013 239 2015 244
rect 2051 252 2053 261
rect 2073 252 2075 261
rect 2084 258 2086 261
rect 2091 258 2093 261
rect 2111 258 2113 261
rect 2121 258 2123 261
rect 2131 266 2133 268
rect 2135 266 2137 268
rect 2131 264 2137 266
rect 2131 251 2133 264
rect 2141 260 2143 273
rect 2158 272 2164 274
rect 2158 270 2160 272
rect 2162 270 2164 272
rect 2158 268 2164 270
rect 2137 258 2143 260
rect 2162 258 2164 268
rect 2169 267 2171 277
rect 2199 285 2205 287
rect 2199 283 2201 285
rect 2203 283 2205 285
rect 2199 281 2208 283
rect 2206 278 2208 281
rect 2182 267 2184 270
rect 2168 265 2174 267
rect 2168 263 2170 265
rect 2172 263 2174 265
rect 2168 261 2174 263
rect 2178 265 2184 267
rect 2178 263 2180 265
rect 2182 263 2184 265
rect 2178 261 2184 263
rect 2172 258 2174 261
rect 2182 258 2184 261
rect 2137 256 2139 258
rect 2141 256 2143 258
rect 2137 254 2143 256
rect 2141 251 2143 254
rect 2111 239 2113 244
rect 2121 239 2123 244
rect 2033 234 2035 238
rect 2040 234 2042 238
rect 2051 234 2053 238
rect 2073 234 2075 238
rect 2084 234 2086 238
rect 2091 234 2093 238
rect 2131 236 2133 241
rect 2162 247 2164 252
rect 2172 247 2174 252
rect 2206 252 2208 270
rect 2216 267 2218 282
rect 2223 277 2225 282
rect 2222 275 2228 277
rect 2222 273 2224 275
rect 2226 273 2228 275
rect 2222 271 2228 273
rect 2233 267 2235 282
rect 2240 272 2242 282
rect 2267 285 2273 287
rect 2267 283 2269 285
rect 2271 283 2273 285
rect 2267 281 2276 283
rect 2212 265 2218 267
rect 2212 263 2214 265
rect 2216 263 2218 265
rect 2212 261 2218 263
rect 2216 252 2218 261
rect 2223 265 2235 267
rect 2239 270 2245 272
rect 2239 268 2241 270
rect 2243 268 2245 270
rect 2239 266 2245 268
rect 2223 252 2225 265
rect 2229 259 2235 261
rect 2229 257 2231 259
rect 2233 257 2235 259
rect 2229 255 2235 257
rect 2233 252 2235 255
rect 2240 252 2242 266
rect 2250 262 2252 280
rect 2274 278 2276 281
rect 2247 260 2253 262
rect 2247 258 2249 260
rect 2251 258 2253 260
rect 2247 256 2253 258
rect 2250 253 2252 256
rect 2182 244 2184 249
rect 2141 234 2143 238
rect 2206 236 2208 246
rect 2274 252 2276 270
rect 2284 267 2286 282
rect 2291 277 2293 282
rect 2290 275 2296 277
rect 2290 273 2292 275
rect 2294 273 2296 275
rect 2290 271 2296 273
rect 2301 267 2303 282
rect 2308 272 2310 282
rect 2280 265 2286 267
rect 2280 263 2282 265
rect 2284 263 2286 265
rect 2280 261 2286 263
rect 2284 252 2286 261
rect 2291 265 2303 267
rect 2307 270 2313 272
rect 2307 268 2309 270
rect 2311 268 2313 270
rect 2307 266 2313 268
rect 2291 252 2293 265
rect 2297 259 2303 261
rect 2297 257 2299 259
rect 2301 257 2303 259
rect 2297 255 2303 257
rect 2301 252 2303 255
rect 2308 252 2310 266
rect 2318 262 2320 280
rect 2315 260 2321 262
rect 2315 258 2317 260
rect 2319 258 2321 260
rect 2315 256 2321 258
rect 2318 253 2320 256
rect 2216 240 2218 244
rect 2223 236 2225 244
rect 2233 239 2235 244
rect 2240 239 2242 244
rect 2250 239 2252 244
rect 2206 234 2225 236
rect 2274 236 2276 246
rect 2284 240 2286 244
rect 2291 236 2293 244
rect 2301 239 2303 244
rect 2308 239 2310 244
rect 2318 239 2320 244
rect 2274 234 2293 236
rect 15 219 17 224
rect 22 219 24 224
rect 35 217 37 221
rect 55 219 57 224
rect 62 219 64 224
rect 95 226 97 230
rect 75 217 77 221
rect 105 223 107 228
rect 145 226 147 230
rect 152 226 154 230
rect 163 226 165 230
rect 185 226 187 230
rect 196 226 198 230
rect 203 226 205 230
rect 115 220 117 225
rect 125 220 127 225
rect 95 210 97 213
rect 95 208 101 210
rect 15 195 17 208
rect 22 203 24 208
rect 35 203 37 208
rect 21 201 27 203
rect 21 199 23 201
rect 25 199 27 201
rect 21 197 27 199
rect 31 201 37 203
rect 31 199 33 201
rect 35 199 37 201
rect 31 197 37 199
rect 11 193 17 195
rect 11 191 13 193
rect 15 191 17 193
rect 11 189 17 191
rect 15 186 17 189
rect 25 186 27 197
rect 35 193 37 197
rect 55 195 57 208
rect 62 203 64 208
rect 75 203 77 208
rect 61 201 67 203
rect 61 199 63 201
rect 65 199 67 201
rect 61 197 67 199
rect 71 201 77 203
rect 71 199 73 201
rect 75 199 77 201
rect 71 197 77 199
rect 51 193 57 195
rect 51 191 53 193
rect 55 191 57 193
rect 51 189 57 191
rect 55 186 57 189
rect 65 186 67 197
rect 75 193 77 197
rect 95 206 97 208
rect 99 206 101 208
rect 95 204 101 206
rect 15 168 17 173
rect 25 168 27 173
rect 35 171 37 175
rect 95 191 97 204
rect 105 200 107 213
rect 101 198 107 200
rect 101 196 103 198
rect 105 196 107 198
rect 115 203 117 206
rect 125 203 127 206
rect 145 203 147 206
rect 152 203 154 206
rect 163 203 165 212
rect 185 203 187 212
rect 223 220 225 225
rect 233 220 235 225
rect 243 223 245 228
rect 253 226 255 230
rect 196 203 198 206
rect 203 203 205 206
rect 223 203 225 206
rect 233 203 235 206
rect 115 201 121 203
rect 115 199 117 201
rect 119 199 121 201
rect 115 197 121 199
rect 125 201 147 203
rect 125 199 136 201
rect 138 199 143 201
rect 145 199 147 201
rect 125 197 147 199
rect 151 201 157 203
rect 151 199 153 201
rect 155 199 157 201
rect 151 197 157 199
rect 161 201 167 203
rect 161 199 163 201
rect 165 199 167 201
rect 161 197 167 199
rect 183 201 189 203
rect 183 199 185 201
rect 187 199 189 201
rect 183 197 189 199
rect 193 201 199 203
rect 193 199 195 201
rect 197 199 199 201
rect 193 197 199 199
rect 203 201 225 203
rect 203 199 205 201
rect 207 199 212 201
rect 214 199 225 201
rect 203 197 225 199
rect 229 201 235 203
rect 229 199 231 201
rect 233 199 235 201
rect 229 197 235 199
rect 243 200 245 213
rect 253 210 255 213
rect 249 208 255 210
rect 249 206 251 208
rect 253 206 255 208
rect 274 212 276 217
rect 284 212 286 217
rect 294 215 296 220
rect 322 219 324 224
rect 329 219 331 224
rect 362 226 364 230
rect 342 217 344 221
rect 372 223 374 228
rect 412 226 414 230
rect 419 226 421 230
rect 430 226 432 230
rect 452 226 454 230
rect 463 226 465 230
rect 470 226 472 230
rect 382 220 384 225
rect 392 220 394 225
rect 362 210 364 213
rect 362 208 368 210
rect 249 204 255 206
rect 243 198 249 200
rect 101 194 110 196
rect 118 194 120 197
rect 125 194 127 197
rect 143 194 145 197
rect 153 194 155 197
rect 163 194 165 197
rect 185 194 187 197
rect 195 194 197 197
rect 205 194 207 197
rect 223 194 225 197
rect 230 194 232 197
rect 243 196 245 198
rect 247 196 249 198
rect 240 194 249 196
rect 108 191 110 194
rect 55 168 57 173
rect 65 168 67 173
rect 75 171 77 175
rect 108 173 110 178
rect 95 162 97 166
rect 118 164 120 169
rect 125 164 127 169
rect 240 191 242 194
rect 253 191 255 204
rect 274 196 276 206
rect 284 203 286 206
rect 294 203 296 206
rect 280 201 286 203
rect 280 199 282 201
rect 284 199 286 201
rect 280 197 286 199
rect 290 201 296 203
rect 290 199 292 201
rect 294 199 296 201
rect 290 197 296 199
rect 270 194 276 196
rect 270 192 272 194
rect 274 192 276 194
rect 240 173 242 178
rect 143 162 145 166
rect 153 162 155 166
rect 163 162 165 166
rect 185 162 187 166
rect 195 162 197 166
rect 205 162 207 166
rect 223 164 225 169
rect 230 164 232 169
rect 270 190 276 192
rect 274 187 276 190
rect 281 187 283 197
rect 294 194 296 197
rect 322 195 324 208
rect 329 203 331 208
rect 342 203 344 208
rect 328 201 334 203
rect 328 199 330 201
rect 332 199 334 201
rect 328 197 334 199
rect 338 201 344 203
rect 338 199 340 201
rect 342 199 344 201
rect 338 197 344 199
rect 318 193 324 195
rect 318 191 320 193
rect 322 191 324 193
rect 318 189 324 191
rect 322 186 324 189
rect 332 186 334 197
rect 342 193 344 197
rect 362 206 364 208
rect 366 206 368 208
rect 362 204 368 206
rect 294 171 296 176
rect 362 191 364 204
rect 372 200 374 213
rect 368 198 374 200
rect 368 196 370 198
rect 372 196 374 198
rect 382 203 384 206
rect 392 203 394 206
rect 412 203 414 206
rect 419 203 421 206
rect 430 203 432 212
rect 452 203 454 212
rect 490 220 492 225
rect 500 220 502 225
rect 510 223 512 228
rect 520 226 522 230
rect 463 203 465 206
rect 470 203 472 206
rect 490 203 492 206
rect 500 203 502 206
rect 382 201 388 203
rect 382 199 384 201
rect 386 199 388 201
rect 382 197 388 199
rect 392 201 414 203
rect 392 199 403 201
rect 405 199 410 201
rect 412 199 414 201
rect 392 197 414 199
rect 418 201 424 203
rect 418 199 420 201
rect 422 199 424 201
rect 418 197 424 199
rect 428 201 434 203
rect 428 199 430 201
rect 432 199 434 201
rect 428 197 434 199
rect 450 201 456 203
rect 450 199 452 201
rect 454 199 456 201
rect 450 197 456 199
rect 460 201 466 203
rect 460 199 462 201
rect 464 199 466 201
rect 460 197 466 199
rect 470 201 492 203
rect 470 199 472 201
rect 474 199 479 201
rect 481 199 492 201
rect 470 197 492 199
rect 496 201 502 203
rect 496 199 498 201
rect 500 199 502 201
rect 496 197 502 199
rect 510 200 512 213
rect 520 210 522 213
rect 516 208 522 210
rect 516 206 518 208
rect 520 206 522 208
rect 541 212 543 217
rect 551 212 553 217
rect 561 215 563 220
rect 589 219 591 224
rect 596 219 598 224
rect 629 226 631 230
rect 609 217 611 221
rect 639 223 641 228
rect 679 226 681 230
rect 686 226 688 230
rect 697 226 699 230
rect 719 226 721 230
rect 730 226 732 230
rect 737 226 739 230
rect 649 220 651 225
rect 659 220 661 225
rect 629 210 631 213
rect 629 208 635 210
rect 516 204 522 206
rect 510 198 516 200
rect 368 194 377 196
rect 385 194 387 197
rect 392 194 394 197
rect 410 194 412 197
rect 420 194 422 197
rect 430 194 432 197
rect 452 194 454 197
rect 462 194 464 197
rect 472 194 474 197
rect 490 194 492 197
rect 497 194 499 197
rect 510 196 512 198
rect 514 196 516 198
rect 507 194 516 196
rect 375 191 377 194
rect 322 168 324 173
rect 332 168 334 173
rect 342 171 344 175
rect 253 162 255 166
rect 274 162 276 166
rect 281 162 283 166
rect 375 173 377 178
rect 362 162 364 166
rect 385 164 387 169
rect 392 164 394 169
rect 507 191 509 194
rect 520 191 522 204
rect 541 196 543 206
rect 551 203 553 206
rect 561 203 563 206
rect 547 201 553 203
rect 547 199 549 201
rect 551 199 553 201
rect 547 197 553 199
rect 557 201 563 203
rect 557 199 559 201
rect 561 199 563 201
rect 557 197 563 199
rect 537 194 543 196
rect 537 192 539 194
rect 541 192 543 194
rect 507 173 509 178
rect 410 162 412 166
rect 420 162 422 166
rect 430 162 432 166
rect 452 162 454 166
rect 462 162 464 166
rect 472 162 474 166
rect 490 164 492 169
rect 497 164 499 169
rect 537 190 543 192
rect 541 187 543 190
rect 548 187 550 197
rect 561 194 563 197
rect 589 195 591 208
rect 596 203 598 208
rect 609 203 611 208
rect 595 201 601 203
rect 595 199 597 201
rect 599 199 601 201
rect 595 197 601 199
rect 605 201 611 203
rect 605 199 607 201
rect 609 199 611 201
rect 605 197 611 199
rect 585 193 591 195
rect 585 191 587 193
rect 589 191 591 193
rect 585 189 591 191
rect 589 186 591 189
rect 599 186 601 197
rect 609 193 611 197
rect 629 206 631 208
rect 633 206 635 208
rect 629 204 635 206
rect 561 171 563 176
rect 629 191 631 204
rect 639 200 641 213
rect 635 198 641 200
rect 635 196 637 198
rect 639 196 641 198
rect 649 203 651 206
rect 659 203 661 206
rect 679 203 681 206
rect 686 203 688 206
rect 697 203 699 212
rect 719 203 721 212
rect 757 220 759 225
rect 767 220 769 225
rect 777 223 779 228
rect 787 226 789 230
rect 730 203 732 206
rect 737 203 739 206
rect 757 203 759 206
rect 767 203 769 206
rect 649 201 655 203
rect 649 199 651 201
rect 653 199 655 201
rect 649 197 655 199
rect 659 201 681 203
rect 659 199 670 201
rect 672 199 677 201
rect 679 199 681 201
rect 659 197 681 199
rect 685 201 691 203
rect 685 199 687 201
rect 689 199 691 201
rect 685 197 691 199
rect 695 201 701 203
rect 695 199 697 201
rect 699 199 701 201
rect 695 197 701 199
rect 717 201 723 203
rect 717 199 719 201
rect 721 199 723 201
rect 717 197 723 199
rect 727 201 733 203
rect 727 199 729 201
rect 731 199 733 201
rect 727 197 733 199
rect 737 201 759 203
rect 737 199 739 201
rect 741 199 746 201
rect 748 199 759 201
rect 737 197 759 199
rect 763 201 769 203
rect 763 199 765 201
rect 767 199 769 201
rect 763 197 769 199
rect 777 200 779 213
rect 787 210 789 213
rect 783 208 789 210
rect 783 206 785 208
rect 787 206 789 208
rect 808 212 810 217
rect 818 212 820 217
rect 828 215 830 220
rect 856 219 858 224
rect 863 219 865 224
rect 896 226 898 230
rect 876 217 878 221
rect 906 223 908 228
rect 946 226 948 230
rect 953 226 955 230
rect 964 226 966 230
rect 986 226 988 230
rect 997 226 999 230
rect 1004 226 1006 230
rect 916 220 918 225
rect 926 220 928 225
rect 896 210 898 213
rect 896 208 902 210
rect 783 204 789 206
rect 777 198 783 200
rect 635 194 644 196
rect 652 194 654 197
rect 659 194 661 197
rect 677 194 679 197
rect 687 194 689 197
rect 697 194 699 197
rect 719 194 721 197
rect 729 194 731 197
rect 739 194 741 197
rect 757 194 759 197
rect 764 194 766 197
rect 777 196 779 198
rect 781 196 783 198
rect 774 194 783 196
rect 642 191 644 194
rect 589 168 591 173
rect 599 168 601 173
rect 609 171 611 175
rect 520 162 522 166
rect 541 162 543 166
rect 548 162 550 166
rect 642 173 644 178
rect 629 162 631 166
rect 652 164 654 169
rect 659 164 661 169
rect 774 191 776 194
rect 787 191 789 204
rect 808 196 810 206
rect 818 203 820 206
rect 828 203 830 206
rect 814 201 820 203
rect 814 199 816 201
rect 818 199 820 201
rect 814 197 820 199
rect 824 201 830 203
rect 824 199 826 201
rect 828 199 830 201
rect 824 197 830 199
rect 804 194 810 196
rect 804 192 806 194
rect 808 192 810 194
rect 774 173 776 178
rect 677 162 679 166
rect 687 162 689 166
rect 697 162 699 166
rect 719 162 721 166
rect 729 162 731 166
rect 739 162 741 166
rect 757 164 759 169
rect 764 164 766 169
rect 804 190 810 192
rect 808 187 810 190
rect 815 187 817 197
rect 828 194 830 197
rect 856 195 858 208
rect 863 203 865 208
rect 876 203 878 208
rect 862 201 868 203
rect 862 199 864 201
rect 866 199 868 201
rect 862 197 868 199
rect 872 201 878 203
rect 872 199 874 201
rect 876 199 878 201
rect 872 197 878 199
rect 852 193 858 195
rect 852 191 854 193
rect 856 191 858 193
rect 852 189 858 191
rect 856 186 858 189
rect 866 186 868 197
rect 876 193 878 197
rect 896 206 898 208
rect 900 206 902 208
rect 896 204 902 206
rect 828 171 830 176
rect 896 191 898 204
rect 906 200 908 213
rect 902 198 908 200
rect 902 196 904 198
rect 906 196 908 198
rect 916 203 918 206
rect 926 203 928 206
rect 946 203 948 206
rect 953 203 955 206
rect 964 203 966 212
rect 986 203 988 212
rect 1024 220 1026 225
rect 1034 220 1036 225
rect 1044 223 1046 228
rect 1054 226 1056 230
rect 997 203 999 206
rect 1004 203 1006 206
rect 1024 203 1026 206
rect 1034 203 1036 206
rect 916 201 922 203
rect 916 199 918 201
rect 920 199 922 201
rect 916 197 922 199
rect 926 201 948 203
rect 926 199 937 201
rect 939 199 944 201
rect 946 199 948 201
rect 926 197 948 199
rect 952 201 958 203
rect 952 199 954 201
rect 956 199 958 201
rect 952 197 958 199
rect 962 201 968 203
rect 962 199 964 201
rect 966 199 968 201
rect 962 197 968 199
rect 984 201 990 203
rect 984 199 986 201
rect 988 199 990 201
rect 984 197 990 199
rect 994 201 1000 203
rect 994 199 996 201
rect 998 199 1000 201
rect 994 197 1000 199
rect 1004 201 1026 203
rect 1004 199 1006 201
rect 1008 199 1013 201
rect 1015 199 1026 201
rect 1004 197 1026 199
rect 1030 201 1036 203
rect 1030 199 1032 201
rect 1034 199 1036 201
rect 1030 197 1036 199
rect 1044 200 1046 213
rect 1054 210 1056 213
rect 1050 208 1056 210
rect 1050 206 1052 208
rect 1054 206 1056 208
rect 1075 212 1077 217
rect 1085 212 1087 217
rect 1095 215 1097 220
rect 1123 219 1125 224
rect 1130 219 1132 224
rect 1163 226 1165 230
rect 1143 217 1145 221
rect 1173 223 1175 228
rect 1213 226 1215 230
rect 1220 226 1222 230
rect 1231 226 1233 230
rect 1253 226 1255 230
rect 1264 226 1266 230
rect 1271 226 1273 230
rect 1183 220 1185 225
rect 1193 220 1195 225
rect 1163 210 1165 213
rect 1163 208 1169 210
rect 1050 204 1056 206
rect 1044 198 1050 200
rect 902 194 911 196
rect 919 194 921 197
rect 926 194 928 197
rect 944 194 946 197
rect 954 194 956 197
rect 964 194 966 197
rect 986 194 988 197
rect 996 194 998 197
rect 1006 194 1008 197
rect 1024 194 1026 197
rect 1031 194 1033 197
rect 1044 196 1046 198
rect 1048 196 1050 198
rect 1041 194 1050 196
rect 909 191 911 194
rect 856 168 858 173
rect 866 168 868 173
rect 876 171 878 175
rect 787 162 789 166
rect 808 162 810 166
rect 815 162 817 166
rect 909 173 911 178
rect 896 162 898 166
rect 919 164 921 169
rect 926 164 928 169
rect 1041 191 1043 194
rect 1054 191 1056 204
rect 1075 196 1077 206
rect 1085 203 1087 206
rect 1095 203 1097 206
rect 1081 201 1087 203
rect 1081 199 1083 201
rect 1085 199 1087 201
rect 1081 197 1087 199
rect 1091 201 1097 203
rect 1091 199 1093 201
rect 1095 199 1097 201
rect 1091 197 1097 199
rect 1071 194 1077 196
rect 1071 192 1073 194
rect 1075 192 1077 194
rect 1041 173 1043 178
rect 944 162 946 166
rect 954 162 956 166
rect 964 162 966 166
rect 986 162 988 166
rect 996 162 998 166
rect 1006 162 1008 166
rect 1024 164 1026 169
rect 1031 164 1033 169
rect 1071 190 1077 192
rect 1075 187 1077 190
rect 1082 187 1084 197
rect 1095 194 1097 197
rect 1123 195 1125 208
rect 1130 203 1132 208
rect 1143 203 1145 208
rect 1129 201 1135 203
rect 1129 199 1131 201
rect 1133 199 1135 201
rect 1129 197 1135 199
rect 1139 201 1145 203
rect 1139 199 1141 201
rect 1143 199 1145 201
rect 1139 197 1145 199
rect 1119 193 1125 195
rect 1119 191 1121 193
rect 1123 191 1125 193
rect 1119 189 1125 191
rect 1123 186 1125 189
rect 1133 186 1135 197
rect 1143 193 1145 197
rect 1163 206 1165 208
rect 1167 206 1169 208
rect 1163 204 1169 206
rect 1095 171 1097 176
rect 1163 191 1165 204
rect 1173 200 1175 213
rect 1169 198 1175 200
rect 1169 196 1171 198
rect 1173 196 1175 198
rect 1183 203 1185 206
rect 1193 203 1195 206
rect 1213 203 1215 206
rect 1220 203 1222 206
rect 1231 203 1233 212
rect 1253 203 1255 212
rect 1291 220 1293 225
rect 1301 220 1303 225
rect 1311 223 1313 228
rect 1321 226 1323 230
rect 1264 203 1266 206
rect 1271 203 1273 206
rect 1291 203 1293 206
rect 1301 203 1303 206
rect 1183 201 1189 203
rect 1183 199 1185 201
rect 1187 199 1189 201
rect 1183 197 1189 199
rect 1193 201 1215 203
rect 1193 199 1204 201
rect 1206 199 1211 201
rect 1213 199 1215 201
rect 1193 197 1215 199
rect 1219 201 1225 203
rect 1219 199 1221 201
rect 1223 199 1225 201
rect 1219 197 1225 199
rect 1229 201 1235 203
rect 1229 199 1231 201
rect 1233 199 1235 201
rect 1229 197 1235 199
rect 1251 201 1257 203
rect 1251 199 1253 201
rect 1255 199 1257 201
rect 1251 197 1257 199
rect 1261 201 1267 203
rect 1261 199 1263 201
rect 1265 199 1267 201
rect 1261 197 1267 199
rect 1271 201 1293 203
rect 1271 199 1273 201
rect 1275 199 1280 201
rect 1282 199 1293 201
rect 1271 197 1293 199
rect 1297 201 1303 203
rect 1297 199 1299 201
rect 1301 199 1303 201
rect 1297 197 1303 199
rect 1311 200 1313 213
rect 1321 210 1323 213
rect 1317 208 1323 210
rect 1317 206 1319 208
rect 1321 206 1323 208
rect 1342 212 1344 217
rect 1352 212 1354 217
rect 1362 215 1364 220
rect 1390 219 1392 224
rect 1397 219 1399 224
rect 1430 226 1432 230
rect 1410 217 1412 221
rect 1440 223 1442 228
rect 1480 226 1482 230
rect 1487 226 1489 230
rect 1498 226 1500 230
rect 1520 226 1522 230
rect 1531 226 1533 230
rect 1538 226 1540 230
rect 1450 220 1452 225
rect 1460 220 1462 225
rect 1430 210 1432 213
rect 1430 208 1436 210
rect 1317 204 1323 206
rect 1311 198 1317 200
rect 1169 194 1178 196
rect 1186 194 1188 197
rect 1193 194 1195 197
rect 1211 194 1213 197
rect 1221 194 1223 197
rect 1231 194 1233 197
rect 1253 194 1255 197
rect 1263 194 1265 197
rect 1273 194 1275 197
rect 1291 194 1293 197
rect 1298 194 1300 197
rect 1311 196 1313 198
rect 1315 196 1317 198
rect 1308 194 1317 196
rect 1176 191 1178 194
rect 1123 168 1125 173
rect 1133 168 1135 173
rect 1143 171 1145 175
rect 1054 162 1056 166
rect 1075 162 1077 166
rect 1082 162 1084 166
rect 1176 173 1178 178
rect 1163 162 1165 166
rect 1186 164 1188 169
rect 1193 164 1195 169
rect 1308 191 1310 194
rect 1321 191 1323 204
rect 1342 196 1344 206
rect 1352 203 1354 206
rect 1362 203 1364 206
rect 1348 201 1354 203
rect 1348 199 1350 201
rect 1352 199 1354 201
rect 1348 197 1354 199
rect 1358 201 1364 203
rect 1358 199 1360 201
rect 1362 199 1364 201
rect 1358 197 1364 199
rect 1338 194 1344 196
rect 1338 192 1340 194
rect 1342 192 1344 194
rect 1308 173 1310 178
rect 1211 162 1213 166
rect 1221 162 1223 166
rect 1231 162 1233 166
rect 1253 162 1255 166
rect 1263 162 1265 166
rect 1273 162 1275 166
rect 1291 164 1293 169
rect 1298 164 1300 169
rect 1338 190 1344 192
rect 1342 187 1344 190
rect 1349 187 1351 197
rect 1362 194 1364 197
rect 1390 195 1392 208
rect 1397 203 1399 208
rect 1410 203 1412 208
rect 1396 201 1402 203
rect 1396 199 1398 201
rect 1400 199 1402 201
rect 1396 197 1402 199
rect 1406 201 1412 203
rect 1406 199 1408 201
rect 1410 199 1412 201
rect 1406 197 1412 199
rect 1386 193 1392 195
rect 1386 191 1388 193
rect 1390 191 1392 193
rect 1386 189 1392 191
rect 1390 186 1392 189
rect 1400 186 1402 197
rect 1410 193 1412 197
rect 1430 206 1432 208
rect 1434 206 1436 208
rect 1430 204 1436 206
rect 1362 171 1364 176
rect 1430 191 1432 204
rect 1440 200 1442 213
rect 1436 198 1442 200
rect 1436 196 1438 198
rect 1440 196 1442 198
rect 1450 203 1452 206
rect 1460 203 1462 206
rect 1480 203 1482 206
rect 1487 203 1489 206
rect 1498 203 1500 212
rect 1520 203 1522 212
rect 1558 220 1560 225
rect 1568 220 1570 225
rect 1578 223 1580 228
rect 1588 226 1590 230
rect 1531 203 1533 206
rect 1538 203 1540 206
rect 1558 203 1560 206
rect 1568 203 1570 206
rect 1450 201 1456 203
rect 1450 199 1452 201
rect 1454 199 1456 201
rect 1450 197 1456 199
rect 1460 201 1482 203
rect 1460 199 1471 201
rect 1473 199 1478 201
rect 1480 199 1482 201
rect 1460 197 1482 199
rect 1486 201 1492 203
rect 1486 199 1488 201
rect 1490 199 1492 201
rect 1486 197 1492 199
rect 1496 201 1502 203
rect 1496 199 1498 201
rect 1500 199 1502 201
rect 1496 197 1502 199
rect 1518 201 1524 203
rect 1518 199 1520 201
rect 1522 199 1524 201
rect 1518 197 1524 199
rect 1528 201 1534 203
rect 1528 199 1530 201
rect 1532 199 1534 201
rect 1528 197 1534 199
rect 1538 201 1560 203
rect 1538 199 1540 201
rect 1542 199 1547 201
rect 1549 199 1560 201
rect 1538 197 1560 199
rect 1564 201 1570 203
rect 1564 199 1566 201
rect 1568 199 1570 201
rect 1564 197 1570 199
rect 1578 200 1580 213
rect 1588 210 1590 213
rect 1584 208 1590 210
rect 1584 206 1586 208
rect 1588 206 1590 208
rect 1609 212 1611 217
rect 1619 212 1621 217
rect 1629 215 1631 220
rect 1657 219 1659 224
rect 1664 219 1666 224
rect 1697 226 1699 230
rect 1677 217 1679 221
rect 1707 223 1709 228
rect 1747 226 1749 230
rect 1754 226 1756 230
rect 1765 226 1767 230
rect 1787 226 1789 230
rect 1798 226 1800 230
rect 1805 226 1807 230
rect 1717 220 1719 225
rect 1727 220 1729 225
rect 1697 210 1699 213
rect 1697 208 1703 210
rect 1584 204 1590 206
rect 1578 198 1584 200
rect 1436 194 1445 196
rect 1453 194 1455 197
rect 1460 194 1462 197
rect 1478 194 1480 197
rect 1488 194 1490 197
rect 1498 194 1500 197
rect 1520 194 1522 197
rect 1530 194 1532 197
rect 1540 194 1542 197
rect 1558 194 1560 197
rect 1565 194 1567 197
rect 1578 196 1580 198
rect 1582 196 1584 198
rect 1575 194 1584 196
rect 1443 191 1445 194
rect 1390 168 1392 173
rect 1400 168 1402 173
rect 1410 171 1412 175
rect 1321 162 1323 166
rect 1342 162 1344 166
rect 1349 162 1351 166
rect 1443 173 1445 178
rect 1430 162 1432 166
rect 1453 164 1455 169
rect 1460 164 1462 169
rect 1575 191 1577 194
rect 1588 191 1590 204
rect 1609 196 1611 206
rect 1619 203 1621 206
rect 1629 203 1631 206
rect 1615 201 1621 203
rect 1615 199 1617 201
rect 1619 199 1621 201
rect 1615 197 1621 199
rect 1625 201 1631 203
rect 1625 199 1627 201
rect 1629 199 1631 201
rect 1625 197 1631 199
rect 1605 194 1611 196
rect 1605 192 1607 194
rect 1609 192 1611 194
rect 1575 173 1577 178
rect 1478 162 1480 166
rect 1488 162 1490 166
rect 1498 162 1500 166
rect 1520 162 1522 166
rect 1530 162 1532 166
rect 1540 162 1542 166
rect 1558 164 1560 169
rect 1565 164 1567 169
rect 1605 190 1611 192
rect 1609 187 1611 190
rect 1616 187 1618 197
rect 1629 194 1631 197
rect 1657 195 1659 208
rect 1664 203 1666 208
rect 1677 203 1679 208
rect 1663 201 1669 203
rect 1663 199 1665 201
rect 1667 199 1669 201
rect 1663 197 1669 199
rect 1673 201 1679 203
rect 1673 199 1675 201
rect 1677 199 1679 201
rect 1673 197 1679 199
rect 1653 193 1659 195
rect 1653 191 1655 193
rect 1657 191 1659 193
rect 1653 189 1659 191
rect 1657 186 1659 189
rect 1667 186 1669 197
rect 1677 193 1679 197
rect 1697 206 1699 208
rect 1701 206 1703 208
rect 1697 204 1703 206
rect 1629 171 1631 176
rect 1697 191 1699 204
rect 1707 200 1709 213
rect 1703 198 1709 200
rect 1703 196 1705 198
rect 1707 196 1709 198
rect 1717 203 1719 206
rect 1727 203 1729 206
rect 1747 203 1749 206
rect 1754 203 1756 206
rect 1765 203 1767 212
rect 1787 203 1789 212
rect 1825 220 1827 225
rect 1835 220 1837 225
rect 1845 223 1847 228
rect 1855 226 1857 230
rect 1922 228 1947 230
rect 1922 220 1924 228
rect 1935 220 1937 224
rect 1945 220 1947 228
rect 1955 223 1957 228
rect 1962 223 1964 228
rect 1983 226 1985 230
rect 1798 203 1800 206
rect 1805 203 1807 206
rect 1825 203 1827 206
rect 1835 203 1837 206
rect 1717 201 1723 203
rect 1717 199 1719 201
rect 1721 199 1723 201
rect 1717 197 1723 199
rect 1727 201 1749 203
rect 1727 199 1738 201
rect 1740 199 1745 201
rect 1747 199 1749 201
rect 1727 197 1749 199
rect 1753 201 1759 203
rect 1753 199 1755 201
rect 1757 199 1759 201
rect 1753 197 1759 199
rect 1763 201 1769 203
rect 1763 199 1765 201
rect 1767 199 1769 201
rect 1763 197 1769 199
rect 1785 201 1791 203
rect 1785 199 1787 201
rect 1789 199 1791 201
rect 1785 197 1791 199
rect 1795 201 1801 203
rect 1795 199 1797 201
rect 1799 199 1801 201
rect 1795 197 1801 199
rect 1805 201 1827 203
rect 1805 199 1807 201
rect 1809 199 1814 201
rect 1816 199 1827 201
rect 1805 197 1827 199
rect 1831 201 1837 203
rect 1831 199 1833 201
rect 1835 199 1837 201
rect 1831 197 1837 199
rect 1845 200 1847 213
rect 1855 210 1857 213
rect 1851 208 1857 210
rect 1851 206 1853 208
rect 1855 206 1857 208
rect 1876 212 1878 217
rect 1886 212 1888 217
rect 1896 215 1898 220
rect 1919 218 1924 220
rect 1919 215 1921 218
rect 1993 223 1995 228
rect 2033 226 2035 230
rect 2040 226 2042 230
rect 2051 226 2053 230
rect 2073 226 2075 230
rect 2084 226 2086 230
rect 2091 226 2093 230
rect 2003 220 2005 225
rect 2013 220 2015 225
rect 1935 208 1937 211
rect 1928 206 1937 208
rect 1945 207 1947 211
rect 1955 208 1957 211
rect 1851 204 1857 206
rect 1845 198 1851 200
rect 1703 194 1712 196
rect 1720 194 1722 197
rect 1727 194 1729 197
rect 1745 194 1747 197
rect 1755 194 1757 197
rect 1765 194 1767 197
rect 1787 194 1789 197
rect 1797 194 1799 197
rect 1807 194 1809 197
rect 1825 194 1827 197
rect 1832 194 1834 197
rect 1845 196 1847 198
rect 1849 196 1851 198
rect 1842 194 1851 196
rect 1710 191 1712 194
rect 1657 168 1659 173
rect 1667 168 1669 173
rect 1677 171 1679 175
rect 1588 162 1590 166
rect 1609 162 1611 166
rect 1616 162 1618 166
rect 1710 173 1712 178
rect 1697 162 1699 166
rect 1720 164 1722 169
rect 1727 164 1729 169
rect 1842 191 1844 194
rect 1855 191 1857 204
rect 1876 196 1878 206
rect 1886 203 1888 206
rect 1896 203 1898 206
rect 1882 201 1888 203
rect 1882 199 1884 201
rect 1886 199 1888 201
rect 1882 197 1888 199
rect 1892 201 1898 203
rect 1892 199 1894 201
rect 1896 199 1898 201
rect 1892 197 1898 199
rect 1919 198 1921 206
rect 1928 204 1930 206
rect 1932 204 1937 206
rect 1928 202 1937 204
rect 1953 206 1957 208
rect 1953 203 1955 206
rect 1935 198 1937 202
rect 1949 201 1955 203
rect 1962 202 1964 211
rect 1983 210 1985 213
rect 1983 208 1989 210
rect 1983 206 1985 208
rect 1987 206 1989 208
rect 1983 204 1989 206
rect 1949 199 1951 201
rect 1953 199 1955 201
rect 1872 194 1878 196
rect 1872 192 1874 194
rect 1876 192 1878 194
rect 1842 173 1844 178
rect 1745 162 1747 166
rect 1755 162 1757 166
rect 1765 162 1767 166
rect 1787 162 1789 166
rect 1797 162 1799 166
rect 1807 162 1809 166
rect 1825 164 1827 169
rect 1832 164 1834 169
rect 1872 190 1878 192
rect 1876 187 1878 190
rect 1883 187 1885 197
rect 1896 194 1898 197
rect 1916 196 1929 198
rect 1935 196 1945 198
rect 1949 197 1955 199
rect 1916 195 1918 196
rect 1912 193 1918 195
rect 1927 193 1929 196
rect 1943 193 1945 196
rect 1953 193 1955 197
rect 1959 200 1965 202
rect 1959 198 1961 200
rect 1963 198 1965 200
rect 1959 196 1965 198
rect 1963 193 1965 196
rect 1912 191 1914 193
rect 1916 191 1918 193
rect 1912 189 1918 191
rect 1896 171 1898 176
rect 1855 162 1857 166
rect 1876 162 1878 166
rect 1883 162 1885 166
rect 1943 171 1945 175
rect 1953 171 1955 175
rect 1927 162 1929 166
rect 1983 191 1985 204
rect 1993 200 1995 213
rect 1989 198 1995 200
rect 1989 196 1991 198
rect 1993 196 1995 198
rect 2003 203 2005 206
rect 2013 203 2015 206
rect 2033 203 2035 206
rect 2040 203 2042 206
rect 2051 203 2053 212
rect 2073 203 2075 212
rect 2111 220 2113 225
rect 2121 220 2123 225
rect 2131 223 2133 228
rect 2141 226 2143 230
rect 2206 228 2225 230
rect 2084 203 2086 206
rect 2091 203 2093 206
rect 2111 203 2113 206
rect 2121 203 2123 206
rect 2003 201 2009 203
rect 2003 199 2005 201
rect 2007 199 2009 201
rect 2003 197 2009 199
rect 2013 201 2035 203
rect 2013 199 2024 201
rect 2026 199 2031 201
rect 2033 199 2035 201
rect 2013 197 2035 199
rect 2039 201 2045 203
rect 2039 199 2041 201
rect 2043 199 2045 201
rect 2039 197 2045 199
rect 2049 201 2055 203
rect 2049 199 2051 201
rect 2053 199 2055 201
rect 2049 197 2055 199
rect 2071 201 2077 203
rect 2071 199 2073 201
rect 2075 199 2077 201
rect 2071 197 2077 199
rect 2081 201 2087 203
rect 2081 199 2083 201
rect 2085 199 2087 201
rect 2081 197 2087 199
rect 2091 201 2113 203
rect 2091 199 2093 201
rect 2095 199 2100 201
rect 2102 199 2113 201
rect 2091 197 2113 199
rect 2117 201 2123 203
rect 2117 199 2119 201
rect 2121 199 2123 201
rect 2117 197 2123 199
rect 2131 200 2133 213
rect 2141 210 2143 213
rect 2137 208 2143 210
rect 2137 206 2139 208
rect 2141 206 2143 208
rect 2162 212 2164 217
rect 2172 212 2174 217
rect 2182 215 2184 220
rect 2206 218 2208 228
rect 2216 220 2218 224
rect 2223 220 2225 228
rect 2274 228 2293 230
rect 2233 220 2235 225
rect 2240 220 2242 225
rect 2250 220 2252 225
rect 2137 204 2143 206
rect 2131 198 2137 200
rect 1989 194 1998 196
rect 2006 194 2008 197
rect 2013 194 2015 197
rect 2031 194 2033 197
rect 2041 194 2043 197
rect 2051 194 2053 197
rect 2073 194 2075 197
rect 2083 194 2085 197
rect 2093 194 2095 197
rect 2111 194 2113 197
rect 2118 194 2120 197
rect 2131 196 2133 198
rect 2135 196 2137 198
rect 2128 194 2137 196
rect 1996 191 1998 194
rect 1996 173 1998 178
rect 1963 162 1965 166
rect 1983 162 1985 166
rect 2006 164 2008 169
rect 2013 164 2015 169
rect 2128 191 2130 194
rect 2141 191 2143 204
rect 2162 196 2164 206
rect 2172 203 2174 206
rect 2182 203 2184 206
rect 2168 201 2174 203
rect 2168 199 2170 201
rect 2172 199 2174 201
rect 2168 197 2174 199
rect 2178 201 2184 203
rect 2178 199 2180 201
rect 2182 199 2184 201
rect 2178 197 2184 199
rect 2158 194 2164 196
rect 2158 192 2160 194
rect 2162 192 2164 194
rect 2128 173 2130 178
rect 2031 162 2033 166
rect 2041 162 2043 166
rect 2051 162 2053 166
rect 2073 162 2075 166
rect 2083 162 2085 166
rect 2093 162 2095 166
rect 2111 164 2113 169
rect 2118 164 2120 169
rect 2158 190 2164 192
rect 2162 187 2164 190
rect 2169 187 2171 197
rect 2182 194 2184 197
rect 2206 194 2208 212
rect 2216 203 2218 212
rect 2212 201 2218 203
rect 2212 199 2214 201
rect 2216 199 2218 201
rect 2212 197 2218 199
rect 2223 199 2225 212
rect 2233 209 2235 212
rect 2229 207 2235 209
rect 2229 205 2231 207
rect 2233 205 2235 207
rect 2229 203 2235 205
rect 2223 197 2235 199
rect 2240 198 2242 212
rect 2274 218 2276 228
rect 2284 220 2286 224
rect 2291 220 2293 228
rect 2301 220 2303 225
rect 2308 220 2310 225
rect 2318 220 2320 225
rect 2250 208 2252 211
rect 2247 206 2253 208
rect 2247 204 2249 206
rect 2251 204 2253 206
rect 2247 202 2253 204
rect 2206 183 2208 186
rect 2199 181 2208 183
rect 2216 182 2218 197
rect 2222 191 2228 193
rect 2222 189 2224 191
rect 2226 189 2228 191
rect 2222 187 2228 189
rect 2223 182 2225 187
rect 2233 182 2235 197
rect 2239 196 2245 198
rect 2239 194 2241 196
rect 2243 194 2245 196
rect 2239 192 2245 194
rect 2240 182 2242 192
rect 2250 184 2252 202
rect 2274 194 2276 212
rect 2284 203 2286 212
rect 2280 201 2286 203
rect 2280 199 2282 201
rect 2284 199 2286 201
rect 2280 197 2286 199
rect 2291 199 2293 212
rect 2301 209 2303 212
rect 2297 207 2303 209
rect 2297 205 2299 207
rect 2301 205 2303 207
rect 2297 203 2303 205
rect 2291 197 2303 199
rect 2308 198 2310 212
rect 2318 208 2320 211
rect 2315 206 2321 208
rect 2315 204 2317 206
rect 2319 204 2321 206
rect 2315 202 2321 204
rect 2199 179 2201 181
rect 2203 179 2205 181
rect 2199 177 2205 179
rect 2182 171 2184 176
rect 2141 162 2143 166
rect 2162 162 2164 166
rect 2169 162 2171 166
rect 2274 183 2276 186
rect 2267 181 2276 183
rect 2284 182 2286 197
rect 2290 191 2296 193
rect 2290 189 2292 191
rect 2294 189 2296 191
rect 2290 187 2296 189
rect 2291 182 2293 187
rect 2301 182 2303 197
rect 2307 196 2313 198
rect 2307 194 2309 196
rect 2311 194 2313 196
rect 2307 192 2313 194
rect 2308 182 2310 192
rect 2318 184 2320 202
rect 2267 179 2269 181
rect 2271 179 2273 181
rect 2267 177 2273 179
rect 2216 162 2218 166
rect 2223 162 2225 166
rect 2233 162 2235 166
rect 2240 162 2242 166
rect 2250 162 2252 166
rect 2284 162 2286 166
rect 2291 162 2293 166
rect 2301 162 2303 166
rect 2308 162 2310 166
rect 2318 162 2320 166
rect 15 147 17 152
rect 25 147 27 152
rect 95 154 97 158
rect 35 145 37 149
rect 55 147 57 152
rect 65 147 67 152
rect 15 131 17 134
rect 11 129 17 131
rect 11 127 13 129
rect 15 127 17 129
rect 11 125 17 127
rect 15 112 17 125
rect 25 123 27 134
rect 75 145 77 149
rect 55 131 57 134
rect 51 129 57 131
rect 51 127 53 129
rect 55 127 57 129
rect 35 123 37 127
rect 51 125 57 127
rect 21 121 27 123
rect 21 119 23 121
rect 25 119 27 121
rect 21 117 27 119
rect 31 121 37 123
rect 31 119 33 121
rect 35 119 37 121
rect 31 117 37 119
rect 22 112 24 117
rect 35 112 37 117
rect 55 112 57 125
rect 65 123 67 134
rect 118 151 120 156
rect 125 151 127 156
rect 143 154 145 158
rect 153 154 155 158
rect 163 154 165 158
rect 185 154 187 158
rect 195 154 197 158
rect 205 154 207 158
rect 108 142 110 147
rect 75 123 77 127
rect 61 121 67 123
rect 61 119 63 121
rect 65 119 67 121
rect 61 117 67 119
rect 71 121 77 123
rect 71 119 73 121
rect 75 119 77 121
rect 71 117 77 119
rect 62 112 64 117
rect 75 112 77 117
rect 95 116 97 129
rect 108 126 110 129
rect 223 151 225 156
rect 230 151 232 156
rect 253 154 255 158
rect 274 154 276 158
rect 281 154 283 158
rect 240 142 242 147
rect 362 154 364 158
rect 294 144 296 149
rect 322 147 324 152
rect 332 147 334 152
rect 274 130 276 133
rect 240 126 242 129
rect 101 124 110 126
rect 101 122 103 124
rect 105 122 107 124
rect 118 123 120 126
rect 125 123 127 126
rect 143 123 145 126
rect 153 123 155 126
rect 163 123 165 126
rect 185 123 187 126
rect 195 123 197 126
rect 205 123 207 126
rect 223 123 225 126
rect 230 123 232 126
rect 240 124 249 126
rect 101 120 107 122
rect 95 114 101 116
rect 95 112 97 114
rect 99 112 101 114
rect 15 96 17 101
rect 22 96 24 101
rect 35 99 37 103
rect 95 110 101 112
rect 95 107 97 110
rect 105 107 107 120
rect 115 121 121 123
rect 115 119 117 121
rect 119 119 121 121
rect 115 117 121 119
rect 125 121 147 123
rect 125 119 136 121
rect 138 119 143 121
rect 145 119 147 121
rect 125 117 147 119
rect 151 121 157 123
rect 151 119 153 121
rect 155 119 157 121
rect 151 117 157 119
rect 161 121 167 123
rect 161 119 163 121
rect 165 119 167 121
rect 161 117 167 119
rect 183 121 189 123
rect 183 119 185 121
rect 187 119 189 121
rect 183 117 189 119
rect 193 121 199 123
rect 193 119 195 121
rect 197 119 199 121
rect 193 117 199 119
rect 203 121 225 123
rect 203 119 205 121
rect 207 119 212 121
rect 214 119 225 121
rect 203 117 225 119
rect 229 121 235 123
rect 229 119 231 121
rect 233 119 235 121
rect 229 117 235 119
rect 115 114 117 117
rect 125 114 127 117
rect 145 114 147 117
rect 152 114 154 117
rect 55 96 57 101
rect 62 96 64 101
rect 75 99 77 103
rect 95 90 97 94
rect 105 92 107 97
rect 115 95 117 100
rect 125 95 127 100
rect 163 108 165 117
rect 185 108 187 117
rect 196 114 198 117
rect 203 114 205 117
rect 223 114 225 117
rect 233 114 235 117
rect 243 122 245 124
rect 247 122 249 124
rect 243 120 249 122
rect 243 107 245 120
rect 253 116 255 129
rect 270 128 276 130
rect 270 126 272 128
rect 274 126 276 128
rect 270 124 276 126
rect 249 114 255 116
rect 274 114 276 124
rect 281 123 283 133
rect 342 145 344 149
rect 322 131 324 134
rect 318 129 324 131
rect 318 127 320 129
rect 322 127 324 129
rect 294 123 296 126
rect 318 125 324 127
rect 280 121 286 123
rect 280 119 282 121
rect 284 119 286 121
rect 280 117 286 119
rect 290 121 296 123
rect 290 119 292 121
rect 294 119 296 121
rect 290 117 296 119
rect 284 114 286 117
rect 294 114 296 117
rect 249 112 251 114
rect 253 112 255 114
rect 249 110 255 112
rect 253 107 255 110
rect 223 95 225 100
rect 233 95 235 100
rect 145 90 147 94
rect 152 90 154 94
rect 163 90 165 94
rect 185 90 187 94
rect 196 90 198 94
rect 203 90 205 94
rect 243 92 245 97
rect 274 103 276 108
rect 284 103 286 108
rect 322 112 324 125
rect 332 123 334 134
rect 385 151 387 156
rect 392 151 394 156
rect 410 154 412 158
rect 420 154 422 158
rect 430 154 432 158
rect 452 154 454 158
rect 462 154 464 158
rect 472 154 474 158
rect 375 142 377 147
rect 342 123 344 127
rect 328 121 334 123
rect 328 119 330 121
rect 332 119 334 121
rect 328 117 334 119
rect 338 121 344 123
rect 338 119 340 121
rect 342 119 344 121
rect 338 117 344 119
rect 329 112 331 117
rect 342 112 344 117
rect 362 116 364 129
rect 375 126 377 129
rect 490 151 492 156
rect 497 151 499 156
rect 520 154 522 158
rect 541 154 543 158
rect 548 154 550 158
rect 507 142 509 147
rect 629 154 631 158
rect 561 144 563 149
rect 589 147 591 152
rect 599 147 601 152
rect 541 130 543 133
rect 507 126 509 129
rect 368 124 377 126
rect 368 122 370 124
rect 372 122 374 124
rect 385 123 387 126
rect 392 123 394 126
rect 410 123 412 126
rect 420 123 422 126
rect 430 123 432 126
rect 452 123 454 126
rect 462 123 464 126
rect 472 123 474 126
rect 490 123 492 126
rect 497 123 499 126
rect 507 124 516 126
rect 368 120 374 122
rect 362 114 368 116
rect 362 112 364 114
rect 366 112 368 114
rect 294 100 296 105
rect 362 110 368 112
rect 362 107 364 110
rect 372 107 374 120
rect 382 121 388 123
rect 382 119 384 121
rect 386 119 388 121
rect 382 117 388 119
rect 392 121 414 123
rect 392 119 403 121
rect 405 119 410 121
rect 412 119 414 121
rect 392 117 414 119
rect 418 121 424 123
rect 418 119 420 121
rect 422 119 424 121
rect 418 117 424 119
rect 428 121 434 123
rect 428 119 430 121
rect 432 119 434 121
rect 428 117 434 119
rect 450 121 456 123
rect 450 119 452 121
rect 454 119 456 121
rect 450 117 456 119
rect 460 121 466 123
rect 460 119 462 121
rect 464 119 466 121
rect 460 117 466 119
rect 470 121 492 123
rect 470 119 472 121
rect 474 119 479 121
rect 481 119 492 121
rect 470 117 492 119
rect 496 121 502 123
rect 496 119 498 121
rect 500 119 502 121
rect 496 117 502 119
rect 382 114 384 117
rect 392 114 394 117
rect 412 114 414 117
rect 419 114 421 117
rect 322 96 324 101
rect 329 96 331 101
rect 253 90 255 94
rect 342 99 344 103
rect 362 90 364 94
rect 372 92 374 97
rect 382 95 384 100
rect 392 95 394 100
rect 430 108 432 117
rect 452 108 454 117
rect 463 114 465 117
rect 470 114 472 117
rect 490 114 492 117
rect 500 114 502 117
rect 510 122 512 124
rect 514 122 516 124
rect 510 120 516 122
rect 510 107 512 120
rect 520 116 522 129
rect 537 128 543 130
rect 537 126 539 128
rect 541 126 543 128
rect 537 124 543 126
rect 516 114 522 116
rect 541 114 543 124
rect 548 123 550 133
rect 609 145 611 149
rect 589 131 591 134
rect 585 129 591 131
rect 585 127 587 129
rect 589 127 591 129
rect 561 123 563 126
rect 585 125 591 127
rect 547 121 553 123
rect 547 119 549 121
rect 551 119 553 121
rect 547 117 553 119
rect 557 121 563 123
rect 557 119 559 121
rect 561 119 563 121
rect 557 117 563 119
rect 551 114 553 117
rect 561 114 563 117
rect 516 112 518 114
rect 520 112 522 114
rect 516 110 522 112
rect 520 107 522 110
rect 490 95 492 100
rect 500 95 502 100
rect 412 90 414 94
rect 419 90 421 94
rect 430 90 432 94
rect 452 90 454 94
rect 463 90 465 94
rect 470 90 472 94
rect 510 92 512 97
rect 541 103 543 108
rect 551 103 553 108
rect 589 112 591 125
rect 599 123 601 134
rect 652 151 654 156
rect 659 151 661 156
rect 677 154 679 158
rect 687 154 689 158
rect 697 154 699 158
rect 719 154 721 158
rect 729 154 731 158
rect 739 154 741 158
rect 642 142 644 147
rect 609 123 611 127
rect 595 121 601 123
rect 595 119 597 121
rect 599 119 601 121
rect 595 117 601 119
rect 605 121 611 123
rect 605 119 607 121
rect 609 119 611 121
rect 605 117 611 119
rect 596 112 598 117
rect 609 112 611 117
rect 629 116 631 129
rect 642 126 644 129
rect 757 151 759 156
rect 764 151 766 156
rect 787 154 789 158
rect 808 154 810 158
rect 815 154 817 158
rect 774 142 776 147
rect 896 154 898 158
rect 828 144 830 149
rect 856 147 858 152
rect 866 147 868 152
rect 808 130 810 133
rect 774 126 776 129
rect 635 124 644 126
rect 635 122 637 124
rect 639 122 641 124
rect 652 123 654 126
rect 659 123 661 126
rect 677 123 679 126
rect 687 123 689 126
rect 697 123 699 126
rect 719 123 721 126
rect 729 123 731 126
rect 739 123 741 126
rect 757 123 759 126
rect 764 123 766 126
rect 774 124 783 126
rect 635 120 641 122
rect 629 114 635 116
rect 629 112 631 114
rect 633 112 635 114
rect 561 100 563 105
rect 629 110 635 112
rect 629 107 631 110
rect 639 107 641 120
rect 649 121 655 123
rect 649 119 651 121
rect 653 119 655 121
rect 649 117 655 119
rect 659 121 681 123
rect 659 119 670 121
rect 672 119 677 121
rect 679 119 681 121
rect 659 117 681 119
rect 685 121 691 123
rect 685 119 687 121
rect 689 119 691 121
rect 685 117 691 119
rect 695 121 701 123
rect 695 119 697 121
rect 699 119 701 121
rect 695 117 701 119
rect 717 121 723 123
rect 717 119 719 121
rect 721 119 723 121
rect 717 117 723 119
rect 727 121 733 123
rect 727 119 729 121
rect 731 119 733 121
rect 727 117 733 119
rect 737 121 759 123
rect 737 119 739 121
rect 741 119 746 121
rect 748 119 759 121
rect 737 117 759 119
rect 763 121 769 123
rect 763 119 765 121
rect 767 119 769 121
rect 763 117 769 119
rect 649 114 651 117
rect 659 114 661 117
rect 679 114 681 117
rect 686 114 688 117
rect 589 96 591 101
rect 596 96 598 101
rect 520 90 522 94
rect 609 99 611 103
rect 629 90 631 94
rect 639 92 641 97
rect 649 95 651 100
rect 659 95 661 100
rect 697 108 699 117
rect 719 108 721 117
rect 730 114 732 117
rect 737 114 739 117
rect 757 114 759 117
rect 767 114 769 117
rect 777 122 779 124
rect 781 122 783 124
rect 777 120 783 122
rect 777 107 779 120
rect 787 116 789 129
rect 804 128 810 130
rect 804 126 806 128
rect 808 126 810 128
rect 804 124 810 126
rect 783 114 789 116
rect 808 114 810 124
rect 815 123 817 133
rect 876 145 878 149
rect 856 131 858 134
rect 852 129 858 131
rect 852 127 854 129
rect 856 127 858 129
rect 828 123 830 126
rect 852 125 858 127
rect 814 121 820 123
rect 814 119 816 121
rect 818 119 820 121
rect 814 117 820 119
rect 824 121 830 123
rect 824 119 826 121
rect 828 119 830 121
rect 824 117 830 119
rect 818 114 820 117
rect 828 114 830 117
rect 783 112 785 114
rect 787 112 789 114
rect 783 110 789 112
rect 787 107 789 110
rect 757 95 759 100
rect 767 95 769 100
rect 679 90 681 94
rect 686 90 688 94
rect 697 90 699 94
rect 719 90 721 94
rect 730 90 732 94
rect 737 90 739 94
rect 777 92 779 97
rect 808 103 810 108
rect 818 103 820 108
rect 856 112 858 125
rect 866 123 868 134
rect 919 151 921 156
rect 926 151 928 156
rect 944 154 946 158
rect 954 154 956 158
rect 964 154 966 158
rect 986 154 988 158
rect 996 154 998 158
rect 1006 154 1008 158
rect 909 142 911 147
rect 876 123 878 127
rect 862 121 868 123
rect 862 119 864 121
rect 866 119 868 121
rect 862 117 868 119
rect 872 121 878 123
rect 872 119 874 121
rect 876 119 878 121
rect 872 117 878 119
rect 863 112 865 117
rect 876 112 878 117
rect 896 116 898 129
rect 909 126 911 129
rect 1024 151 1026 156
rect 1031 151 1033 156
rect 1054 154 1056 158
rect 1075 154 1077 158
rect 1082 154 1084 158
rect 1041 142 1043 147
rect 1163 154 1165 158
rect 1095 144 1097 149
rect 1123 147 1125 152
rect 1133 147 1135 152
rect 1075 130 1077 133
rect 1041 126 1043 129
rect 902 124 911 126
rect 902 122 904 124
rect 906 122 908 124
rect 919 123 921 126
rect 926 123 928 126
rect 944 123 946 126
rect 954 123 956 126
rect 964 123 966 126
rect 986 123 988 126
rect 996 123 998 126
rect 1006 123 1008 126
rect 1024 123 1026 126
rect 1031 123 1033 126
rect 1041 124 1050 126
rect 902 120 908 122
rect 896 114 902 116
rect 896 112 898 114
rect 900 112 902 114
rect 828 100 830 105
rect 896 110 902 112
rect 896 107 898 110
rect 906 107 908 120
rect 916 121 922 123
rect 916 119 918 121
rect 920 119 922 121
rect 916 117 922 119
rect 926 121 948 123
rect 926 119 937 121
rect 939 119 944 121
rect 946 119 948 121
rect 926 117 948 119
rect 952 121 958 123
rect 952 119 954 121
rect 956 119 958 121
rect 952 117 958 119
rect 962 121 968 123
rect 962 119 964 121
rect 966 119 968 121
rect 962 117 968 119
rect 984 121 990 123
rect 984 119 986 121
rect 988 119 990 121
rect 984 117 990 119
rect 994 121 1000 123
rect 994 119 996 121
rect 998 119 1000 121
rect 994 117 1000 119
rect 1004 121 1026 123
rect 1004 119 1006 121
rect 1008 119 1013 121
rect 1015 119 1026 121
rect 1004 117 1026 119
rect 1030 121 1036 123
rect 1030 119 1032 121
rect 1034 119 1036 121
rect 1030 117 1036 119
rect 916 114 918 117
rect 926 114 928 117
rect 946 114 948 117
rect 953 114 955 117
rect 856 96 858 101
rect 863 96 865 101
rect 787 90 789 94
rect 876 99 878 103
rect 896 90 898 94
rect 906 92 908 97
rect 916 95 918 100
rect 926 95 928 100
rect 964 108 966 117
rect 986 108 988 117
rect 997 114 999 117
rect 1004 114 1006 117
rect 1024 114 1026 117
rect 1034 114 1036 117
rect 1044 122 1046 124
rect 1048 122 1050 124
rect 1044 120 1050 122
rect 1044 107 1046 120
rect 1054 116 1056 129
rect 1071 128 1077 130
rect 1071 126 1073 128
rect 1075 126 1077 128
rect 1071 124 1077 126
rect 1050 114 1056 116
rect 1075 114 1077 124
rect 1082 123 1084 133
rect 1143 145 1145 149
rect 1123 131 1125 134
rect 1119 129 1125 131
rect 1119 127 1121 129
rect 1123 127 1125 129
rect 1095 123 1097 126
rect 1119 125 1125 127
rect 1081 121 1087 123
rect 1081 119 1083 121
rect 1085 119 1087 121
rect 1081 117 1087 119
rect 1091 121 1097 123
rect 1091 119 1093 121
rect 1095 119 1097 121
rect 1091 117 1097 119
rect 1085 114 1087 117
rect 1095 114 1097 117
rect 1050 112 1052 114
rect 1054 112 1056 114
rect 1050 110 1056 112
rect 1054 107 1056 110
rect 1024 95 1026 100
rect 1034 95 1036 100
rect 946 90 948 94
rect 953 90 955 94
rect 964 90 966 94
rect 986 90 988 94
rect 997 90 999 94
rect 1004 90 1006 94
rect 1044 92 1046 97
rect 1075 103 1077 108
rect 1085 103 1087 108
rect 1123 112 1125 125
rect 1133 123 1135 134
rect 1186 151 1188 156
rect 1193 151 1195 156
rect 1211 154 1213 158
rect 1221 154 1223 158
rect 1231 154 1233 158
rect 1253 154 1255 158
rect 1263 154 1265 158
rect 1273 154 1275 158
rect 1176 142 1178 147
rect 1143 123 1145 127
rect 1129 121 1135 123
rect 1129 119 1131 121
rect 1133 119 1135 121
rect 1129 117 1135 119
rect 1139 121 1145 123
rect 1139 119 1141 121
rect 1143 119 1145 121
rect 1139 117 1145 119
rect 1130 112 1132 117
rect 1143 112 1145 117
rect 1163 116 1165 129
rect 1176 126 1178 129
rect 1291 151 1293 156
rect 1298 151 1300 156
rect 1321 154 1323 158
rect 1342 154 1344 158
rect 1349 154 1351 158
rect 1308 142 1310 147
rect 1430 154 1432 158
rect 1362 144 1364 149
rect 1390 147 1392 152
rect 1400 147 1402 152
rect 1342 130 1344 133
rect 1308 126 1310 129
rect 1169 124 1178 126
rect 1169 122 1171 124
rect 1173 122 1175 124
rect 1186 123 1188 126
rect 1193 123 1195 126
rect 1211 123 1213 126
rect 1221 123 1223 126
rect 1231 123 1233 126
rect 1253 123 1255 126
rect 1263 123 1265 126
rect 1273 123 1275 126
rect 1291 123 1293 126
rect 1298 123 1300 126
rect 1308 124 1317 126
rect 1169 120 1175 122
rect 1163 114 1169 116
rect 1163 112 1165 114
rect 1167 112 1169 114
rect 1095 100 1097 105
rect 1163 110 1169 112
rect 1163 107 1165 110
rect 1173 107 1175 120
rect 1183 121 1189 123
rect 1183 119 1185 121
rect 1187 119 1189 121
rect 1183 117 1189 119
rect 1193 121 1215 123
rect 1193 119 1204 121
rect 1206 119 1211 121
rect 1213 119 1215 121
rect 1193 117 1215 119
rect 1219 121 1225 123
rect 1219 119 1221 121
rect 1223 119 1225 121
rect 1219 117 1225 119
rect 1229 121 1235 123
rect 1229 119 1231 121
rect 1233 119 1235 121
rect 1229 117 1235 119
rect 1251 121 1257 123
rect 1251 119 1253 121
rect 1255 119 1257 121
rect 1251 117 1257 119
rect 1261 121 1267 123
rect 1261 119 1263 121
rect 1265 119 1267 121
rect 1261 117 1267 119
rect 1271 121 1293 123
rect 1271 119 1273 121
rect 1275 119 1280 121
rect 1282 119 1293 121
rect 1271 117 1293 119
rect 1297 121 1303 123
rect 1297 119 1299 121
rect 1301 119 1303 121
rect 1297 117 1303 119
rect 1183 114 1185 117
rect 1193 114 1195 117
rect 1213 114 1215 117
rect 1220 114 1222 117
rect 1123 96 1125 101
rect 1130 96 1132 101
rect 1054 90 1056 94
rect 1143 99 1145 103
rect 1163 90 1165 94
rect 1173 92 1175 97
rect 1183 95 1185 100
rect 1193 95 1195 100
rect 1231 108 1233 117
rect 1253 108 1255 117
rect 1264 114 1266 117
rect 1271 114 1273 117
rect 1291 114 1293 117
rect 1301 114 1303 117
rect 1311 122 1313 124
rect 1315 122 1317 124
rect 1311 120 1317 122
rect 1311 107 1313 120
rect 1321 116 1323 129
rect 1338 128 1344 130
rect 1338 126 1340 128
rect 1342 126 1344 128
rect 1338 124 1344 126
rect 1317 114 1323 116
rect 1342 114 1344 124
rect 1349 123 1351 133
rect 1410 145 1412 149
rect 1390 131 1392 134
rect 1386 129 1392 131
rect 1386 127 1388 129
rect 1390 127 1392 129
rect 1362 123 1364 126
rect 1386 125 1392 127
rect 1348 121 1354 123
rect 1348 119 1350 121
rect 1352 119 1354 121
rect 1348 117 1354 119
rect 1358 121 1364 123
rect 1358 119 1360 121
rect 1362 119 1364 121
rect 1358 117 1364 119
rect 1352 114 1354 117
rect 1362 114 1364 117
rect 1317 112 1319 114
rect 1321 112 1323 114
rect 1317 110 1323 112
rect 1321 107 1323 110
rect 1291 95 1293 100
rect 1301 95 1303 100
rect 1213 90 1215 94
rect 1220 90 1222 94
rect 1231 90 1233 94
rect 1253 90 1255 94
rect 1264 90 1266 94
rect 1271 90 1273 94
rect 1311 92 1313 97
rect 1342 103 1344 108
rect 1352 103 1354 108
rect 1390 112 1392 125
rect 1400 123 1402 134
rect 1453 151 1455 156
rect 1460 151 1462 156
rect 1478 154 1480 158
rect 1488 154 1490 158
rect 1498 154 1500 158
rect 1520 154 1522 158
rect 1530 154 1532 158
rect 1540 154 1542 158
rect 1443 142 1445 147
rect 1410 123 1412 127
rect 1396 121 1402 123
rect 1396 119 1398 121
rect 1400 119 1402 121
rect 1396 117 1402 119
rect 1406 121 1412 123
rect 1406 119 1408 121
rect 1410 119 1412 121
rect 1406 117 1412 119
rect 1397 112 1399 117
rect 1410 112 1412 117
rect 1430 116 1432 129
rect 1443 126 1445 129
rect 1558 151 1560 156
rect 1565 151 1567 156
rect 1588 154 1590 158
rect 1609 154 1611 158
rect 1616 154 1618 158
rect 1575 142 1577 147
rect 1697 154 1699 158
rect 1629 144 1631 149
rect 1657 147 1659 152
rect 1667 147 1669 152
rect 1609 130 1611 133
rect 1575 126 1577 129
rect 1436 124 1445 126
rect 1436 122 1438 124
rect 1440 122 1442 124
rect 1453 123 1455 126
rect 1460 123 1462 126
rect 1478 123 1480 126
rect 1488 123 1490 126
rect 1498 123 1500 126
rect 1520 123 1522 126
rect 1530 123 1532 126
rect 1540 123 1542 126
rect 1558 123 1560 126
rect 1565 123 1567 126
rect 1575 124 1584 126
rect 1436 120 1442 122
rect 1430 114 1436 116
rect 1430 112 1432 114
rect 1434 112 1436 114
rect 1362 100 1364 105
rect 1430 110 1436 112
rect 1430 107 1432 110
rect 1440 107 1442 120
rect 1450 121 1456 123
rect 1450 119 1452 121
rect 1454 119 1456 121
rect 1450 117 1456 119
rect 1460 121 1482 123
rect 1460 119 1471 121
rect 1473 119 1478 121
rect 1480 119 1482 121
rect 1460 117 1482 119
rect 1486 121 1492 123
rect 1486 119 1488 121
rect 1490 119 1492 121
rect 1486 117 1492 119
rect 1496 121 1502 123
rect 1496 119 1498 121
rect 1500 119 1502 121
rect 1496 117 1502 119
rect 1518 121 1524 123
rect 1518 119 1520 121
rect 1522 119 1524 121
rect 1518 117 1524 119
rect 1528 121 1534 123
rect 1528 119 1530 121
rect 1532 119 1534 121
rect 1528 117 1534 119
rect 1538 121 1560 123
rect 1538 119 1540 121
rect 1542 119 1547 121
rect 1549 119 1560 121
rect 1538 117 1560 119
rect 1564 121 1570 123
rect 1564 119 1566 121
rect 1568 119 1570 121
rect 1564 117 1570 119
rect 1450 114 1452 117
rect 1460 114 1462 117
rect 1480 114 1482 117
rect 1487 114 1489 117
rect 1390 96 1392 101
rect 1397 96 1399 101
rect 1321 90 1323 94
rect 1410 99 1412 103
rect 1430 90 1432 94
rect 1440 92 1442 97
rect 1450 95 1452 100
rect 1460 95 1462 100
rect 1498 108 1500 117
rect 1520 108 1522 117
rect 1531 114 1533 117
rect 1538 114 1540 117
rect 1558 114 1560 117
rect 1568 114 1570 117
rect 1578 122 1580 124
rect 1582 122 1584 124
rect 1578 120 1584 122
rect 1578 107 1580 120
rect 1588 116 1590 129
rect 1605 128 1611 130
rect 1605 126 1607 128
rect 1609 126 1611 128
rect 1605 124 1611 126
rect 1584 114 1590 116
rect 1609 114 1611 124
rect 1616 123 1618 133
rect 1677 145 1679 149
rect 1657 131 1659 134
rect 1653 129 1659 131
rect 1653 127 1655 129
rect 1657 127 1659 129
rect 1629 123 1631 126
rect 1653 125 1659 127
rect 1615 121 1621 123
rect 1615 119 1617 121
rect 1619 119 1621 121
rect 1615 117 1621 119
rect 1625 121 1631 123
rect 1625 119 1627 121
rect 1629 119 1631 121
rect 1625 117 1631 119
rect 1619 114 1621 117
rect 1629 114 1631 117
rect 1584 112 1586 114
rect 1588 112 1590 114
rect 1584 110 1590 112
rect 1588 107 1590 110
rect 1558 95 1560 100
rect 1568 95 1570 100
rect 1480 90 1482 94
rect 1487 90 1489 94
rect 1498 90 1500 94
rect 1520 90 1522 94
rect 1531 90 1533 94
rect 1538 90 1540 94
rect 1578 92 1580 97
rect 1609 103 1611 108
rect 1619 103 1621 108
rect 1657 112 1659 125
rect 1667 123 1669 134
rect 1720 151 1722 156
rect 1727 151 1729 156
rect 1745 154 1747 158
rect 1755 154 1757 158
rect 1765 154 1767 158
rect 1787 154 1789 158
rect 1797 154 1799 158
rect 1807 154 1809 158
rect 1710 142 1712 147
rect 1677 123 1679 127
rect 1663 121 1669 123
rect 1663 119 1665 121
rect 1667 119 1669 121
rect 1663 117 1669 119
rect 1673 121 1679 123
rect 1673 119 1675 121
rect 1677 119 1679 121
rect 1673 117 1679 119
rect 1664 112 1666 117
rect 1677 112 1679 117
rect 1697 116 1699 129
rect 1710 126 1712 129
rect 1825 151 1827 156
rect 1832 151 1834 156
rect 1855 154 1857 158
rect 1876 154 1878 158
rect 1883 154 1885 158
rect 1842 142 1844 147
rect 1927 154 1929 158
rect 1896 144 1898 149
rect 1876 130 1878 133
rect 1842 126 1844 129
rect 1703 124 1712 126
rect 1703 122 1705 124
rect 1707 122 1709 124
rect 1720 123 1722 126
rect 1727 123 1729 126
rect 1745 123 1747 126
rect 1755 123 1757 126
rect 1765 123 1767 126
rect 1787 123 1789 126
rect 1797 123 1799 126
rect 1807 123 1809 126
rect 1825 123 1827 126
rect 1832 123 1834 126
rect 1842 124 1851 126
rect 1703 120 1709 122
rect 1697 114 1703 116
rect 1697 112 1699 114
rect 1701 112 1703 114
rect 1629 100 1631 105
rect 1697 110 1703 112
rect 1697 107 1699 110
rect 1707 107 1709 120
rect 1717 121 1723 123
rect 1717 119 1719 121
rect 1721 119 1723 121
rect 1717 117 1723 119
rect 1727 121 1749 123
rect 1727 119 1738 121
rect 1740 119 1745 121
rect 1747 119 1749 121
rect 1727 117 1749 119
rect 1753 121 1759 123
rect 1753 119 1755 121
rect 1757 119 1759 121
rect 1753 117 1759 119
rect 1763 121 1769 123
rect 1763 119 1765 121
rect 1767 119 1769 121
rect 1763 117 1769 119
rect 1785 121 1791 123
rect 1785 119 1787 121
rect 1789 119 1791 121
rect 1785 117 1791 119
rect 1795 121 1801 123
rect 1795 119 1797 121
rect 1799 119 1801 121
rect 1795 117 1801 119
rect 1805 121 1827 123
rect 1805 119 1807 121
rect 1809 119 1814 121
rect 1816 119 1827 121
rect 1805 117 1827 119
rect 1831 121 1837 123
rect 1831 119 1833 121
rect 1835 119 1837 121
rect 1831 117 1837 119
rect 1717 114 1719 117
rect 1727 114 1729 117
rect 1747 114 1749 117
rect 1754 114 1756 117
rect 1657 96 1659 101
rect 1664 96 1666 101
rect 1588 90 1590 94
rect 1677 99 1679 103
rect 1697 90 1699 94
rect 1707 92 1709 97
rect 1717 95 1719 100
rect 1727 95 1729 100
rect 1765 108 1767 117
rect 1787 108 1789 117
rect 1798 114 1800 117
rect 1805 114 1807 117
rect 1825 114 1827 117
rect 1835 114 1837 117
rect 1845 122 1847 124
rect 1849 122 1851 124
rect 1845 120 1851 122
rect 1845 107 1847 120
rect 1855 116 1857 129
rect 1872 128 1878 130
rect 1872 126 1874 128
rect 1876 126 1878 128
rect 1872 124 1878 126
rect 1851 114 1857 116
rect 1876 114 1878 124
rect 1883 123 1885 133
rect 1912 129 1918 131
rect 1912 127 1914 129
rect 1916 127 1918 129
rect 1963 154 1965 158
rect 1983 154 1985 158
rect 1943 145 1945 149
rect 1953 145 1955 149
rect 2006 151 2008 156
rect 2013 151 2015 156
rect 2031 154 2033 158
rect 2041 154 2043 158
rect 2051 154 2053 158
rect 2073 154 2075 158
rect 2083 154 2085 158
rect 2093 154 2095 158
rect 1996 142 1998 147
rect 1896 123 1898 126
rect 1912 125 1918 127
rect 1882 121 1888 123
rect 1882 119 1884 121
rect 1886 119 1888 121
rect 1882 117 1888 119
rect 1892 121 1898 123
rect 1916 124 1918 125
rect 1927 124 1929 127
rect 1943 124 1945 127
rect 1916 122 1929 124
rect 1935 122 1945 124
rect 1953 123 1955 127
rect 1963 124 1965 127
rect 1892 119 1894 121
rect 1896 119 1898 121
rect 1892 117 1898 119
rect 1886 114 1888 117
rect 1896 114 1898 117
rect 1919 114 1921 122
rect 1935 118 1937 122
rect 1928 116 1937 118
rect 1949 121 1955 123
rect 1949 119 1951 121
rect 1953 119 1955 121
rect 1949 117 1955 119
rect 1959 122 1965 124
rect 1959 120 1961 122
rect 1963 120 1965 122
rect 1959 118 1965 120
rect 1928 114 1930 116
rect 1932 114 1937 116
rect 1851 112 1853 114
rect 1855 112 1857 114
rect 1851 110 1857 112
rect 1855 107 1857 110
rect 1825 95 1827 100
rect 1835 95 1837 100
rect 1747 90 1749 94
rect 1754 90 1756 94
rect 1765 90 1767 94
rect 1787 90 1789 94
rect 1798 90 1800 94
rect 1805 90 1807 94
rect 1845 92 1847 97
rect 1876 103 1878 108
rect 1886 103 1888 108
rect 1928 112 1937 114
rect 1953 114 1955 117
rect 1935 109 1937 112
rect 1945 109 1947 113
rect 1953 112 1957 114
rect 1955 109 1957 112
rect 1962 109 1964 118
rect 1983 116 1985 129
rect 1996 126 1998 129
rect 2111 151 2113 156
rect 2118 151 2120 156
rect 2141 154 2143 158
rect 2162 154 2164 158
rect 2169 154 2171 158
rect 2128 142 2130 147
rect 2216 154 2218 158
rect 2223 154 2225 158
rect 2233 154 2235 158
rect 2240 154 2242 158
rect 2250 154 2252 158
rect 2284 154 2286 158
rect 2291 154 2293 158
rect 2301 154 2303 158
rect 2308 154 2310 158
rect 2318 154 2320 158
rect 2182 144 2184 149
rect 2162 130 2164 133
rect 2128 126 2130 129
rect 1989 124 1998 126
rect 1989 122 1991 124
rect 1993 122 1995 124
rect 2006 123 2008 126
rect 2013 123 2015 126
rect 2031 123 2033 126
rect 2041 123 2043 126
rect 2051 123 2053 126
rect 2073 123 2075 126
rect 2083 123 2085 126
rect 2093 123 2095 126
rect 2111 123 2113 126
rect 2118 123 2120 126
rect 2128 124 2137 126
rect 1989 120 1995 122
rect 1983 114 1989 116
rect 1983 112 1985 114
rect 1987 112 1989 114
rect 1983 110 1989 112
rect 1896 100 1898 105
rect 1919 102 1921 105
rect 1919 100 1924 102
rect 1855 90 1857 94
rect 1922 92 1924 100
rect 1935 96 1937 100
rect 1945 92 1947 100
rect 1983 107 1985 110
rect 1993 107 1995 120
rect 2003 121 2009 123
rect 2003 119 2005 121
rect 2007 119 2009 121
rect 2003 117 2009 119
rect 2013 121 2035 123
rect 2013 119 2024 121
rect 2026 119 2031 121
rect 2033 119 2035 121
rect 2013 117 2035 119
rect 2039 121 2045 123
rect 2039 119 2041 121
rect 2043 119 2045 121
rect 2039 117 2045 119
rect 2049 121 2055 123
rect 2049 119 2051 121
rect 2053 119 2055 121
rect 2049 117 2055 119
rect 2071 121 2077 123
rect 2071 119 2073 121
rect 2075 119 2077 121
rect 2071 117 2077 119
rect 2081 121 2087 123
rect 2081 119 2083 121
rect 2085 119 2087 121
rect 2081 117 2087 119
rect 2091 121 2113 123
rect 2091 119 2093 121
rect 2095 119 2100 121
rect 2102 119 2113 121
rect 2091 117 2113 119
rect 2117 121 2123 123
rect 2117 119 2119 121
rect 2121 119 2123 121
rect 2117 117 2123 119
rect 2003 114 2005 117
rect 2013 114 2015 117
rect 2033 114 2035 117
rect 2040 114 2042 117
rect 1955 92 1957 97
rect 1962 92 1964 97
rect 1922 90 1947 92
rect 1983 90 1985 94
rect 1993 92 1995 97
rect 2003 95 2005 100
rect 2013 95 2015 100
rect 2051 108 2053 117
rect 2073 108 2075 117
rect 2084 114 2086 117
rect 2091 114 2093 117
rect 2111 114 2113 117
rect 2121 114 2123 117
rect 2131 122 2133 124
rect 2135 122 2137 124
rect 2131 120 2137 122
rect 2131 107 2133 120
rect 2141 116 2143 129
rect 2158 128 2164 130
rect 2158 126 2160 128
rect 2162 126 2164 128
rect 2158 124 2164 126
rect 2137 114 2143 116
rect 2162 114 2164 124
rect 2169 123 2171 133
rect 2199 141 2205 143
rect 2199 139 2201 141
rect 2203 139 2205 141
rect 2199 137 2208 139
rect 2206 134 2208 137
rect 2182 123 2184 126
rect 2168 121 2174 123
rect 2168 119 2170 121
rect 2172 119 2174 121
rect 2168 117 2174 119
rect 2178 121 2184 123
rect 2178 119 2180 121
rect 2182 119 2184 121
rect 2178 117 2184 119
rect 2172 114 2174 117
rect 2182 114 2184 117
rect 2137 112 2139 114
rect 2141 112 2143 114
rect 2137 110 2143 112
rect 2141 107 2143 110
rect 2111 95 2113 100
rect 2121 95 2123 100
rect 2033 90 2035 94
rect 2040 90 2042 94
rect 2051 90 2053 94
rect 2073 90 2075 94
rect 2084 90 2086 94
rect 2091 90 2093 94
rect 2131 92 2133 97
rect 2162 103 2164 108
rect 2172 103 2174 108
rect 2206 108 2208 126
rect 2216 123 2218 138
rect 2223 133 2225 138
rect 2222 131 2228 133
rect 2222 129 2224 131
rect 2226 129 2228 131
rect 2222 127 2228 129
rect 2233 123 2235 138
rect 2240 128 2242 138
rect 2267 141 2273 143
rect 2267 139 2269 141
rect 2271 139 2273 141
rect 2267 137 2276 139
rect 2212 121 2218 123
rect 2212 119 2214 121
rect 2216 119 2218 121
rect 2212 117 2218 119
rect 2216 108 2218 117
rect 2223 121 2235 123
rect 2239 126 2245 128
rect 2239 124 2241 126
rect 2243 124 2245 126
rect 2239 122 2245 124
rect 2223 108 2225 121
rect 2229 115 2235 117
rect 2229 113 2231 115
rect 2233 113 2235 115
rect 2229 111 2235 113
rect 2233 108 2235 111
rect 2240 108 2242 122
rect 2250 118 2252 136
rect 2274 134 2276 137
rect 2247 116 2253 118
rect 2247 114 2249 116
rect 2251 114 2253 116
rect 2247 112 2253 114
rect 2250 109 2252 112
rect 2182 100 2184 105
rect 2141 90 2143 94
rect 2206 92 2208 102
rect 2274 108 2276 126
rect 2284 123 2286 138
rect 2291 133 2293 138
rect 2290 131 2296 133
rect 2290 129 2292 131
rect 2294 129 2296 131
rect 2290 127 2296 129
rect 2301 123 2303 138
rect 2308 128 2310 138
rect 2280 121 2286 123
rect 2280 119 2282 121
rect 2284 119 2286 121
rect 2280 117 2286 119
rect 2284 108 2286 117
rect 2291 121 2303 123
rect 2307 126 2313 128
rect 2307 124 2309 126
rect 2311 124 2313 126
rect 2307 122 2313 124
rect 2291 108 2293 121
rect 2297 115 2303 117
rect 2297 113 2299 115
rect 2301 113 2303 115
rect 2297 111 2303 113
rect 2301 108 2303 111
rect 2308 108 2310 122
rect 2318 118 2320 136
rect 2315 116 2321 118
rect 2315 114 2317 116
rect 2319 114 2321 116
rect 2315 112 2321 114
rect 2318 109 2320 112
rect 2216 96 2218 100
rect 2223 92 2225 100
rect 2233 95 2235 100
rect 2240 95 2242 100
rect 2250 95 2252 100
rect 2206 90 2225 92
rect 2274 92 2276 102
rect 2284 96 2286 100
rect 2291 92 2293 100
rect 2301 95 2303 100
rect 2308 95 2310 100
rect 2318 95 2320 100
rect 2274 90 2293 92
rect 15 75 17 80
rect 22 75 24 80
rect 35 73 37 77
rect 55 75 57 80
rect 62 75 64 80
rect 95 82 97 86
rect 75 73 77 77
rect 105 79 107 84
rect 145 82 147 86
rect 152 82 154 86
rect 163 82 165 86
rect 185 82 187 86
rect 196 82 198 86
rect 203 82 205 86
rect 115 76 117 81
rect 125 76 127 81
rect 95 66 97 69
rect 95 64 101 66
rect 15 51 17 64
rect 22 59 24 64
rect 35 59 37 64
rect 21 57 27 59
rect 21 55 23 57
rect 25 55 27 57
rect 21 53 27 55
rect 31 57 37 59
rect 31 55 33 57
rect 35 55 37 57
rect 31 53 37 55
rect 11 49 17 51
rect 11 47 13 49
rect 15 47 17 49
rect 11 45 17 47
rect 15 42 17 45
rect 25 42 27 53
rect 35 49 37 53
rect 55 51 57 64
rect 62 59 64 64
rect 75 59 77 64
rect 61 57 67 59
rect 61 55 63 57
rect 65 55 67 57
rect 61 53 67 55
rect 71 57 77 59
rect 71 55 73 57
rect 75 55 77 57
rect 71 53 77 55
rect 51 49 57 51
rect 51 47 53 49
rect 55 47 57 49
rect 51 45 57 47
rect 55 42 57 45
rect 65 42 67 53
rect 75 49 77 53
rect 95 62 97 64
rect 99 62 101 64
rect 95 60 101 62
rect 15 24 17 29
rect 25 24 27 29
rect 35 27 37 31
rect 95 47 97 60
rect 105 56 107 69
rect 101 54 107 56
rect 101 52 103 54
rect 105 52 107 54
rect 115 59 117 62
rect 125 59 127 62
rect 145 59 147 62
rect 152 59 154 62
rect 163 59 165 68
rect 185 59 187 68
rect 223 76 225 81
rect 233 76 235 81
rect 243 79 245 84
rect 253 82 255 86
rect 196 59 198 62
rect 203 59 205 62
rect 223 59 225 62
rect 233 59 235 62
rect 115 57 121 59
rect 115 55 117 57
rect 119 55 121 57
rect 115 53 121 55
rect 125 57 147 59
rect 125 55 136 57
rect 138 55 143 57
rect 145 55 147 57
rect 125 53 147 55
rect 151 57 157 59
rect 151 55 153 57
rect 155 55 157 57
rect 151 53 157 55
rect 161 57 167 59
rect 161 55 163 57
rect 165 55 167 57
rect 161 53 167 55
rect 183 57 189 59
rect 183 55 185 57
rect 187 55 189 57
rect 183 53 189 55
rect 193 57 199 59
rect 193 55 195 57
rect 197 55 199 57
rect 193 53 199 55
rect 203 57 225 59
rect 203 55 205 57
rect 207 55 212 57
rect 214 55 225 57
rect 203 53 225 55
rect 229 57 235 59
rect 229 55 231 57
rect 233 55 235 57
rect 229 53 235 55
rect 243 56 245 69
rect 253 66 255 69
rect 249 64 255 66
rect 249 62 251 64
rect 253 62 255 64
rect 274 68 276 73
rect 284 68 286 73
rect 294 71 296 76
rect 322 75 324 80
rect 329 75 331 80
rect 362 82 364 86
rect 342 73 344 77
rect 372 79 374 84
rect 412 82 414 86
rect 419 82 421 86
rect 430 82 432 86
rect 452 82 454 86
rect 463 82 465 86
rect 470 82 472 86
rect 382 76 384 81
rect 392 76 394 81
rect 362 66 364 69
rect 362 64 368 66
rect 249 60 255 62
rect 243 54 249 56
rect 101 50 110 52
rect 118 50 120 53
rect 125 50 127 53
rect 143 50 145 53
rect 153 50 155 53
rect 163 50 165 53
rect 185 50 187 53
rect 195 50 197 53
rect 205 50 207 53
rect 223 50 225 53
rect 230 50 232 53
rect 243 52 245 54
rect 247 52 249 54
rect 240 50 249 52
rect 108 47 110 50
rect 55 24 57 29
rect 65 24 67 29
rect 75 27 77 31
rect 108 29 110 34
rect 95 18 97 22
rect 118 20 120 25
rect 125 20 127 25
rect 240 47 242 50
rect 253 47 255 60
rect 274 52 276 62
rect 284 59 286 62
rect 294 59 296 62
rect 280 57 286 59
rect 280 55 282 57
rect 284 55 286 57
rect 280 53 286 55
rect 290 57 296 59
rect 290 55 292 57
rect 294 55 296 57
rect 290 53 296 55
rect 270 50 276 52
rect 270 48 272 50
rect 274 48 276 50
rect 240 29 242 34
rect 143 18 145 22
rect 153 18 155 22
rect 163 18 165 22
rect 185 18 187 22
rect 195 18 197 22
rect 205 18 207 22
rect 223 20 225 25
rect 230 20 232 25
rect 270 46 276 48
rect 274 43 276 46
rect 281 43 283 53
rect 294 50 296 53
rect 322 51 324 64
rect 329 59 331 64
rect 342 59 344 64
rect 328 57 334 59
rect 328 55 330 57
rect 332 55 334 57
rect 328 53 334 55
rect 338 57 344 59
rect 338 55 340 57
rect 342 55 344 57
rect 338 53 344 55
rect 318 49 324 51
rect 318 47 320 49
rect 322 47 324 49
rect 318 45 324 47
rect 322 42 324 45
rect 332 42 334 53
rect 342 49 344 53
rect 362 62 364 64
rect 366 62 368 64
rect 362 60 368 62
rect 294 27 296 32
rect 362 47 364 60
rect 372 56 374 69
rect 368 54 374 56
rect 368 52 370 54
rect 372 52 374 54
rect 382 59 384 62
rect 392 59 394 62
rect 412 59 414 62
rect 419 59 421 62
rect 430 59 432 68
rect 452 59 454 68
rect 490 76 492 81
rect 500 76 502 81
rect 510 79 512 84
rect 520 82 522 86
rect 463 59 465 62
rect 470 59 472 62
rect 490 59 492 62
rect 500 59 502 62
rect 382 57 388 59
rect 382 55 384 57
rect 386 55 388 57
rect 382 53 388 55
rect 392 57 414 59
rect 392 55 403 57
rect 405 55 410 57
rect 412 55 414 57
rect 392 53 414 55
rect 418 57 424 59
rect 418 55 420 57
rect 422 55 424 57
rect 418 53 424 55
rect 428 57 434 59
rect 428 55 430 57
rect 432 55 434 57
rect 428 53 434 55
rect 450 57 456 59
rect 450 55 452 57
rect 454 55 456 57
rect 450 53 456 55
rect 460 57 466 59
rect 460 55 462 57
rect 464 55 466 57
rect 460 53 466 55
rect 470 57 492 59
rect 470 55 472 57
rect 474 55 479 57
rect 481 55 492 57
rect 470 53 492 55
rect 496 57 502 59
rect 496 55 498 57
rect 500 55 502 57
rect 496 53 502 55
rect 510 56 512 69
rect 520 66 522 69
rect 516 64 522 66
rect 516 62 518 64
rect 520 62 522 64
rect 541 68 543 73
rect 551 68 553 73
rect 561 71 563 76
rect 589 75 591 80
rect 596 75 598 80
rect 629 82 631 86
rect 609 73 611 77
rect 639 79 641 84
rect 679 82 681 86
rect 686 82 688 86
rect 697 82 699 86
rect 719 82 721 86
rect 730 82 732 86
rect 737 82 739 86
rect 649 76 651 81
rect 659 76 661 81
rect 629 66 631 69
rect 629 64 635 66
rect 516 60 522 62
rect 510 54 516 56
rect 368 50 377 52
rect 385 50 387 53
rect 392 50 394 53
rect 410 50 412 53
rect 420 50 422 53
rect 430 50 432 53
rect 452 50 454 53
rect 462 50 464 53
rect 472 50 474 53
rect 490 50 492 53
rect 497 50 499 53
rect 510 52 512 54
rect 514 52 516 54
rect 507 50 516 52
rect 375 47 377 50
rect 322 24 324 29
rect 332 24 334 29
rect 342 27 344 31
rect 253 18 255 22
rect 274 18 276 22
rect 281 18 283 22
rect 375 29 377 34
rect 362 18 364 22
rect 385 20 387 25
rect 392 20 394 25
rect 507 47 509 50
rect 520 47 522 60
rect 541 52 543 62
rect 551 59 553 62
rect 561 59 563 62
rect 547 57 553 59
rect 547 55 549 57
rect 551 55 553 57
rect 547 53 553 55
rect 557 57 563 59
rect 557 55 559 57
rect 561 55 563 57
rect 557 53 563 55
rect 537 50 543 52
rect 537 48 539 50
rect 541 48 543 50
rect 507 29 509 34
rect 410 18 412 22
rect 420 18 422 22
rect 430 18 432 22
rect 452 18 454 22
rect 462 18 464 22
rect 472 18 474 22
rect 490 20 492 25
rect 497 20 499 25
rect 537 46 543 48
rect 541 43 543 46
rect 548 43 550 53
rect 561 50 563 53
rect 589 51 591 64
rect 596 59 598 64
rect 609 59 611 64
rect 595 57 601 59
rect 595 55 597 57
rect 599 55 601 57
rect 595 53 601 55
rect 605 57 611 59
rect 605 55 607 57
rect 609 55 611 57
rect 605 53 611 55
rect 585 49 591 51
rect 585 47 587 49
rect 589 47 591 49
rect 585 45 591 47
rect 589 42 591 45
rect 599 42 601 53
rect 609 49 611 53
rect 629 62 631 64
rect 633 62 635 64
rect 629 60 635 62
rect 561 27 563 32
rect 629 47 631 60
rect 639 56 641 69
rect 635 54 641 56
rect 635 52 637 54
rect 639 52 641 54
rect 649 59 651 62
rect 659 59 661 62
rect 679 59 681 62
rect 686 59 688 62
rect 697 59 699 68
rect 719 59 721 68
rect 757 76 759 81
rect 767 76 769 81
rect 777 79 779 84
rect 787 82 789 86
rect 730 59 732 62
rect 737 59 739 62
rect 757 59 759 62
rect 767 59 769 62
rect 649 57 655 59
rect 649 55 651 57
rect 653 55 655 57
rect 649 53 655 55
rect 659 57 681 59
rect 659 55 670 57
rect 672 55 677 57
rect 679 55 681 57
rect 659 53 681 55
rect 685 57 691 59
rect 685 55 687 57
rect 689 55 691 57
rect 685 53 691 55
rect 695 57 701 59
rect 695 55 697 57
rect 699 55 701 57
rect 695 53 701 55
rect 717 57 723 59
rect 717 55 719 57
rect 721 55 723 57
rect 717 53 723 55
rect 727 57 733 59
rect 727 55 729 57
rect 731 55 733 57
rect 727 53 733 55
rect 737 57 759 59
rect 737 55 739 57
rect 741 55 746 57
rect 748 55 759 57
rect 737 53 759 55
rect 763 57 769 59
rect 763 55 765 57
rect 767 55 769 57
rect 763 53 769 55
rect 777 56 779 69
rect 787 66 789 69
rect 783 64 789 66
rect 783 62 785 64
rect 787 62 789 64
rect 808 68 810 73
rect 818 68 820 73
rect 828 71 830 76
rect 856 75 858 80
rect 863 75 865 80
rect 896 82 898 86
rect 876 73 878 77
rect 906 79 908 84
rect 946 82 948 86
rect 953 82 955 86
rect 964 82 966 86
rect 986 82 988 86
rect 997 82 999 86
rect 1004 82 1006 86
rect 916 76 918 81
rect 926 76 928 81
rect 896 66 898 69
rect 896 64 902 66
rect 783 60 789 62
rect 777 54 783 56
rect 635 50 644 52
rect 652 50 654 53
rect 659 50 661 53
rect 677 50 679 53
rect 687 50 689 53
rect 697 50 699 53
rect 719 50 721 53
rect 729 50 731 53
rect 739 50 741 53
rect 757 50 759 53
rect 764 50 766 53
rect 777 52 779 54
rect 781 52 783 54
rect 774 50 783 52
rect 642 47 644 50
rect 589 24 591 29
rect 599 24 601 29
rect 609 27 611 31
rect 520 18 522 22
rect 541 18 543 22
rect 548 18 550 22
rect 642 29 644 34
rect 629 18 631 22
rect 652 20 654 25
rect 659 20 661 25
rect 774 47 776 50
rect 787 47 789 60
rect 808 52 810 62
rect 818 59 820 62
rect 828 59 830 62
rect 814 57 820 59
rect 814 55 816 57
rect 818 55 820 57
rect 814 53 820 55
rect 824 57 830 59
rect 824 55 826 57
rect 828 55 830 57
rect 824 53 830 55
rect 804 50 810 52
rect 804 48 806 50
rect 808 48 810 50
rect 774 29 776 34
rect 677 18 679 22
rect 687 18 689 22
rect 697 18 699 22
rect 719 18 721 22
rect 729 18 731 22
rect 739 18 741 22
rect 757 20 759 25
rect 764 20 766 25
rect 804 46 810 48
rect 808 43 810 46
rect 815 43 817 53
rect 828 50 830 53
rect 856 51 858 64
rect 863 59 865 64
rect 876 59 878 64
rect 862 57 868 59
rect 862 55 864 57
rect 866 55 868 57
rect 862 53 868 55
rect 872 57 878 59
rect 872 55 874 57
rect 876 55 878 57
rect 872 53 878 55
rect 852 49 858 51
rect 852 47 854 49
rect 856 47 858 49
rect 852 45 858 47
rect 856 42 858 45
rect 866 42 868 53
rect 876 49 878 53
rect 896 62 898 64
rect 900 62 902 64
rect 896 60 902 62
rect 828 27 830 32
rect 896 47 898 60
rect 906 56 908 69
rect 902 54 908 56
rect 902 52 904 54
rect 906 52 908 54
rect 916 59 918 62
rect 926 59 928 62
rect 946 59 948 62
rect 953 59 955 62
rect 964 59 966 68
rect 986 59 988 68
rect 1024 76 1026 81
rect 1034 76 1036 81
rect 1044 79 1046 84
rect 1054 82 1056 86
rect 997 59 999 62
rect 1004 59 1006 62
rect 1024 59 1026 62
rect 1034 59 1036 62
rect 916 57 922 59
rect 916 55 918 57
rect 920 55 922 57
rect 916 53 922 55
rect 926 57 948 59
rect 926 55 937 57
rect 939 55 944 57
rect 946 55 948 57
rect 926 53 948 55
rect 952 57 958 59
rect 952 55 954 57
rect 956 55 958 57
rect 952 53 958 55
rect 962 57 968 59
rect 962 55 964 57
rect 966 55 968 57
rect 962 53 968 55
rect 984 57 990 59
rect 984 55 986 57
rect 988 55 990 57
rect 984 53 990 55
rect 994 57 1000 59
rect 994 55 996 57
rect 998 55 1000 57
rect 994 53 1000 55
rect 1004 57 1026 59
rect 1004 55 1006 57
rect 1008 55 1013 57
rect 1015 55 1026 57
rect 1004 53 1026 55
rect 1030 57 1036 59
rect 1030 55 1032 57
rect 1034 55 1036 57
rect 1030 53 1036 55
rect 1044 56 1046 69
rect 1054 66 1056 69
rect 1050 64 1056 66
rect 1050 62 1052 64
rect 1054 62 1056 64
rect 1075 68 1077 73
rect 1085 68 1087 73
rect 1095 71 1097 76
rect 1123 75 1125 80
rect 1130 75 1132 80
rect 1163 82 1165 86
rect 1143 73 1145 77
rect 1173 79 1175 84
rect 1213 82 1215 86
rect 1220 82 1222 86
rect 1231 82 1233 86
rect 1253 82 1255 86
rect 1264 82 1266 86
rect 1271 82 1273 86
rect 1183 76 1185 81
rect 1193 76 1195 81
rect 1163 66 1165 69
rect 1163 64 1169 66
rect 1050 60 1056 62
rect 1044 54 1050 56
rect 902 50 911 52
rect 919 50 921 53
rect 926 50 928 53
rect 944 50 946 53
rect 954 50 956 53
rect 964 50 966 53
rect 986 50 988 53
rect 996 50 998 53
rect 1006 50 1008 53
rect 1024 50 1026 53
rect 1031 50 1033 53
rect 1044 52 1046 54
rect 1048 52 1050 54
rect 1041 50 1050 52
rect 909 47 911 50
rect 856 24 858 29
rect 866 24 868 29
rect 876 27 878 31
rect 787 18 789 22
rect 808 18 810 22
rect 815 18 817 22
rect 909 29 911 34
rect 896 18 898 22
rect 919 20 921 25
rect 926 20 928 25
rect 1041 47 1043 50
rect 1054 47 1056 60
rect 1075 52 1077 62
rect 1085 59 1087 62
rect 1095 59 1097 62
rect 1081 57 1087 59
rect 1081 55 1083 57
rect 1085 55 1087 57
rect 1081 53 1087 55
rect 1091 57 1097 59
rect 1091 55 1093 57
rect 1095 55 1097 57
rect 1091 53 1097 55
rect 1071 50 1077 52
rect 1071 48 1073 50
rect 1075 48 1077 50
rect 1041 29 1043 34
rect 944 18 946 22
rect 954 18 956 22
rect 964 18 966 22
rect 986 18 988 22
rect 996 18 998 22
rect 1006 18 1008 22
rect 1024 20 1026 25
rect 1031 20 1033 25
rect 1071 46 1077 48
rect 1075 43 1077 46
rect 1082 43 1084 53
rect 1095 50 1097 53
rect 1123 51 1125 64
rect 1130 59 1132 64
rect 1143 59 1145 64
rect 1129 57 1135 59
rect 1129 55 1131 57
rect 1133 55 1135 57
rect 1129 53 1135 55
rect 1139 57 1145 59
rect 1139 55 1141 57
rect 1143 55 1145 57
rect 1139 53 1145 55
rect 1119 49 1125 51
rect 1119 47 1121 49
rect 1123 47 1125 49
rect 1119 45 1125 47
rect 1123 42 1125 45
rect 1133 42 1135 53
rect 1143 49 1145 53
rect 1163 62 1165 64
rect 1167 62 1169 64
rect 1163 60 1169 62
rect 1095 27 1097 32
rect 1163 47 1165 60
rect 1173 56 1175 69
rect 1169 54 1175 56
rect 1169 52 1171 54
rect 1173 52 1175 54
rect 1183 59 1185 62
rect 1193 59 1195 62
rect 1213 59 1215 62
rect 1220 59 1222 62
rect 1231 59 1233 68
rect 1253 59 1255 68
rect 1291 76 1293 81
rect 1301 76 1303 81
rect 1311 79 1313 84
rect 1321 82 1323 86
rect 1264 59 1266 62
rect 1271 59 1273 62
rect 1291 59 1293 62
rect 1301 59 1303 62
rect 1183 57 1189 59
rect 1183 55 1185 57
rect 1187 55 1189 57
rect 1183 53 1189 55
rect 1193 57 1215 59
rect 1193 55 1204 57
rect 1206 55 1211 57
rect 1213 55 1215 57
rect 1193 53 1215 55
rect 1219 57 1225 59
rect 1219 55 1221 57
rect 1223 55 1225 57
rect 1219 53 1225 55
rect 1229 57 1235 59
rect 1229 55 1231 57
rect 1233 55 1235 57
rect 1229 53 1235 55
rect 1251 57 1257 59
rect 1251 55 1253 57
rect 1255 55 1257 57
rect 1251 53 1257 55
rect 1261 57 1267 59
rect 1261 55 1263 57
rect 1265 55 1267 57
rect 1261 53 1267 55
rect 1271 57 1293 59
rect 1271 55 1273 57
rect 1275 55 1280 57
rect 1282 55 1293 57
rect 1271 53 1293 55
rect 1297 57 1303 59
rect 1297 55 1299 57
rect 1301 55 1303 57
rect 1297 53 1303 55
rect 1311 56 1313 69
rect 1321 66 1323 69
rect 1317 64 1323 66
rect 1317 62 1319 64
rect 1321 62 1323 64
rect 1342 68 1344 73
rect 1352 68 1354 73
rect 1362 71 1364 76
rect 1390 75 1392 80
rect 1397 75 1399 80
rect 1430 82 1432 86
rect 1410 73 1412 77
rect 1440 79 1442 84
rect 1480 82 1482 86
rect 1487 82 1489 86
rect 1498 82 1500 86
rect 1520 82 1522 86
rect 1531 82 1533 86
rect 1538 82 1540 86
rect 1450 76 1452 81
rect 1460 76 1462 81
rect 1430 66 1432 69
rect 1430 64 1436 66
rect 1317 60 1323 62
rect 1311 54 1317 56
rect 1169 50 1178 52
rect 1186 50 1188 53
rect 1193 50 1195 53
rect 1211 50 1213 53
rect 1221 50 1223 53
rect 1231 50 1233 53
rect 1253 50 1255 53
rect 1263 50 1265 53
rect 1273 50 1275 53
rect 1291 50 1293 53
rect 1298 50 1300 53
rect 1311 52 1313 54
rect 1315 52 1317 54
rect 1308 50 1317 52
rect 1176 47 1178 50
rect 1123 24 1125 29
rect 1133 24 1135 29
rect 1143 27 1145 31
rect 1054 18 1056 22
rect 1075 18 1077 22
rect 1082 18 1084 22
rect 1176 29 1178 34
rect 1163 18 1165 22
rect 1186 20 1188 25
rect 1193 20 1195 25
rect 1308 47 1310 50
rect 1321 47 1323 60
rect 1342 52 1344 62
rect 1352 59 1354 62
rect 1362 59 1364 62
rect 1348 57 1354 59
rect 1348 55 1350 57
rect 1352 55 1354 57
rect 1348 53 1354 55
rect 1358 57 1364 59
rect 1358 55 1360 57
rect 1362 55 1364 57
rect 1358 53 1364 55
rect 1338 50 1344 52
rect 1338 48 1340 50
rect 1342 48 1344 50
rect 1308 29 1310 34
rect 1211 18 1213 22
rect 1221 18 1223 22
rect 1231 18 1233 22
rect 1253 18 1255 22
rect 1263 18 1265 22
rect 1273 18 1275 22
rect 1291 20 1293 25
rect 1298 20 1300 25
rect 1338 46 1344 48
rect 1342 43 1344 46
rect 1349 43 1351 53
rect 1362 50 1364 53
rect 1390 51 1392 64
rect 1397 59 1399 64
rect 1410 59 1412 64
rect 1396 57 1402 59
rect 1396 55 1398 57
rect 1400 55 1402 57
rect 1396 53 1402 55
rect 1406 57 1412 59
rect 1406 55 1408 57
rect 1410 55 1412 57
rect 1406 53 1412 55
rect 1386 49 1392 51
rect 1386 47 1388 49
rect 1390 47 1392 49
rect 1386 45 1392 47
rect 1390 42 1392 45
rect 1400 42 1402 53
rect 1410 49 1412 53
rect 1430 62 1432 64
rect 1434 62 1436 64
rect 1430 60 1436 62
rect 1362 27 1364 32
rect 1430 47 1432 60
rect 1440 56 1442 69
rect 1436 54 1442 56
rect 1436 52 1438 54
rect 1440 52 1442 54
rect 1450 59 1452 62
rect 1460 59 1462 62
rect 1480 59 1482 62
rect 1487 59 1489 62
rect 1498 59 1500 68
rect 1520 59 1522 68
rect 1558 76 1560 81
rect 1568 76 1570 81
rect 1578 79 1580 84
rect 1588 82 1590 86
rect 1531 59 1533 62
rect 1538 59 1540 62
rect 1558 59 1560 62
rect 1568 59 1570 62
rect 1450 57 1456 59
rect 1450 55 1452 57
rect 1454 55 1456 57
rect 1450 53 1456 55
rect 1460 57 1482 59
rect 1460 55 1471 57
rect 1473 55 1478 57
rect 1480 55 1482 57
rect 1460 53 1482 55
rect 1486 57 1492 59
rect 1486 55 1488 57
rect 1490 55 1492 57
rect 1486 53 1492 55
rect 1496 57 1502 59
rect 1496 55 1498 57
rect 1500 55 1502 57
rect 1496 53 1502 55
rect 1518 57 1524 59
rect 1518 55 1520 57
rect 1522 55 1524 57
rect 1518 53 1524 55
rect 1528 57 1534 59
rect 1528 55 1530 57
rect 1532 55 1534 57
rect 1528 53 1534 55
rect 1538 57 1560 59
rect 1538 55 1540 57
rect 1542 55 1547 57
rect 1549 55 1560 57
rect 1538 53 1560 55
rect 1564 57 1570 59
rect 1564 55 1566 57
rect 1568 55 1570 57
rect 1564 53 1570 55
rect 1578 56 1580 69
rect 1588 66 1590 69
rect 1584 64 1590 66
rect 1584 62 1586 64
rect 1588 62 1590 64
rect 1609 68 1611 73
rect 1619 68 1621 73
rect 1629 71 1631 76
rect 1657 75 1659 80
rect 1664 75 1666 80
rect 1697 82 1699 86
rect 1677 73 1679 77
rect 1707 79 1709 84
rect 1747 82 1749 86
rect 1754 82 1756 86
rect 1765 82 1767 86
rect 1787 82 1789 86
rect 1798 82 1800 86
rect 1805 82 1807 86
rect 1717 76 1719 81
rect 1727 76 1729 81
rect 1697 66 1699 69
rect 1697 64 1703 66
rect 1584 60 1590 62
rect 1578 54 1584 56
rect 1436 50 1445 52
rect 1453 50 1455 53
rect 1460 50 1462 53
rect 1478 50 1480 53
rect 1488 50 1490 53
rect 1498 50 1500 53
rect 1520 50 1522 53
rect 1530 50 1532 53
rect 1540 50 1542 53
rect 1558 50 1560 53
rect 1565 50 1567 53
rect 1578 52 1580 54
rect 1582 52 1584 54
rect 1575 50 1584 52
rect 1443 47 1445 50
rect 1390 24 1392 29
rect 1400 24 1402 29
rect 1410 27 1412 31
rect 1321 18 1323 22
rect 1342 18 1344 22
rect 1349 18 1351 22
rect 1443 29 1445 34
rect 1430 18 1432 22
rect 1453 20 1455 25
rect 1460 20 1462 25
rect 1575 47 1577 50
rect 1588 47 1590 60
rect 1609 52 1611 62
rect 1619 59 1621 62
rect 1629 59 1631 62
rect 1615 57 1621 59
rect 1615 55 1617 57
rect 1619 55 1621 57
rect 1615 53 1621 55
rect 1625 57 1631 59
rect 1625 55 1627 57
rect 1629 55 1631 57
rect 1625 53 1631 55
rect 1605 50 1611 52
rect 1605 48 1607 50
rect 1609 48 1611 50
rect 1575 29 1577 34
rect 1478 18 1480 22
rect 1488 18 1490 22
rect 1498 18 1500 22
rect 1520 18 1522 22
rect 1530 18 1532 22
rect 1540 18 1542 22
rect 1558 20 1560 25
rect 1565 20 1567 25
rect 1605 46 1611 48
rect 1609 43 1611 46
rect 1616 43 1618 53
rect 1629 50 1631 53
rect 1657 51 1659 64
rect 1664 59 1666 64
rect 1677 59 1679 64
rect 1663 57 1669 59
rect 1663 55 1665 57
rect 1667 55 1669 57
rect 1663 53 1669 55
rect 1673 57 1679 59
rect 1673 55 1675 57
rect 1677 55 1679 57
rect 1673 53 1679 55
rect 1653 49 1659 51
rect 1653 47 1655 49
rect 1657 47 1659 49
rect 1653 45 1659 47
rect 1657 42 1659 45
rect 1667 42 1669 53
rect 1677 49 1679 53
rect 1697 62 1699 64
rect 1701 62 1703 64
rect 1697 60 1703 62
rect 1629 27 1631 32
rect 1697 47 1699 60
rect 1707 56 1709 69
rect 1703 54 1709 56
rect 1703 52 1705 54
rect 1707 52 1709 54
rect 1717 59 1719 62
rect 1727 59 1729 62
rect 1747 59 1749 62
rect 1754 59 1756 62
rect 1765 59 1767 68
rect 1787 59 1789 68
rect 1825 76 1827 81
rect 1835 76 1837 81
rect 1845 79 1847 84
rect 1855 82 1857 86
rect 1922 84 1947 86
rect 1922 76 1924 84
rect 1935 76 1937 80
rect 1945 76 1947 84
rect 1955 79 1957 84
rect 1962 79 1964 84
rect 1983 82 1985 86
rect 1798 59 1800 62
rect 1805 59 1807 62
rect 1825 59 1827 62
rect 1835 59 1837 62
rect 1717 57 1723 59
rect 1717 55 1719 57
rect 1721 55 1723 57
rect 1717 53 1723 55
rect 1727 57 1749 59
rect 1727 55 1738 57
rect 1740 55 1745 57
rect 1747 55 1749 57
rect 1727 53 1749 55
rect 1753 57 1759 59
rect 1753 55 1755 57
rect 1757 55 1759 57
rect 1753 53 1759 55
rect 1763 57 1769 59
rect 1763 55 1765 57
rect 1767 55 1769 57
rect 1763 53 1769 55
rect 1785 57 1791 59
rect 1785 55 1787 57
rect 1789 55 1791 57
rect 1785 53 1791 55
rect 1795 57 1801 59
rect 1795 55 1797 57
rect 1799 55 1801 57
rect 1795 53 1801 55
rect 1805 57 1827 59
rect 1805 55 1807 57
rect 1809 55 1814 57
rect 1816 55 1827 57
rect 1805 53 1827 55
rect 1831 57 1837 59
rect 1831 55 1833 57
rect 1835 55 1837 57
rect 1831 53 1837 55
rect 1845 56 1847 69
rect 1855 66 1857 69
rect 1851 64 1857 66
rect 1851 62 1853 64
rect 1855 62 1857 64
rect 1876 68 1878 73
rect 1886 68 1888 73
rect 1896 71 1898 76
rect 1919 74 1924 76
rect 1919 71 1921 74
rect 1993 79 1995 84
rect 2033 82 2035 86
rect 2040 82 2042 86
rect 2051 82 2053 86
rect 2073 82 2075 86
rect 2084 82 2086 86
rect 2091 82 2093 86
rect 2003 76 2005 81
rect 2013 76 2015 81
rect 1935 64 1937 67
rect 1928 62 1937 64
rect 1945 63 1947 67
rect 1955 64 1957 67
rect 1851 60 1857 62
rect 1845 54 1851 56
rect 1703 50 1712 52
rect 1720 50 1722 53
rect 1727 50 1729 53
rect 1745 50 1747 53
rect 1755 50 1757 53
rect 1765 50 1767 53
rect 1787 50 1789 53
rect 1797 50 1799 53
rect 1807 50 1809 53
rect 1825 50 1827 53
rect 1832 50 1834 53
rect 1845 52 1847 54
rect 1849 52 1851 54
rect 1842 50 1851 52
rect 1710 47 1712 50
rect 1657 24 1659 29
rect 1667 24 1669 29
rect 1677 27 1679 31
rect 1588 18 1590 22
rect 1609 18 1611 22
rect 1616 18 1618 22
rect 1710 29 1712 34
rect 1697 18 1699 22
rect 1720 20 1722 25
rect 1727 20 1729 25
rect 1842 47 1844 50
rect 1855 47 1857 60
rect 1876 52 1878 62
rect 1886 59 1888 62
rect 1896 59 1898 62
rect 1882 57 1888 59
rect 1882 55 1884 57
rect 1886 55 1888 57
rect 1882 53 1888 55
rect 1892 57 1898 59
rect 1892 55 1894 57
rect 1896 55 1898 57
rect 1892 53 1898 55
rect 1919 54 1921 62
rect 1928 60 1930 62
rect 1932 60 1937 62
rect 1928 58 1937 60
rect 1953 62 1957 64
rect 1953 59 1955 62
rect 1935 54 1937 58
rect 1949 57 1955 59
rect 1962 58 1964 67
rect 1983 66 1985 69
rect 1983 64 1989 66
rect 1983 62 1985 64
rect 1987 62 1989 64
rect 1983 60 1989 62
rect 1949 55 1951 57
rect 1953 55 1955 57
rect 1872 50 1878 52
rect 1872 48 1874 50
rect 1876 48 1878 50
rect 1842 29 1844 34
rect 1745 18 1747 22
rect 1755 18 1757 22
rect 1765 18 1767 22
rect 1787 18 1789 22
rect 1797 18 1799 22
rect 1807 18 1809 22
rect 1825 20 1827 25
rect 1832 20 1834 25
rect 1872 46 1878 48
rect 1876 43 1878 46
rect 1883 43 1885 53
rect 1896 50 1898 53
rect 1916 52 1929 54
rect 1935 52 1945 54
rect 1949 53 1955 55
rect 1916 51 1918 52
rect 1912 49 1918 51
rect 1927 49 1929 52
rect 1943 49 1945 52
rect 1953 49 1955 53
rect 1959 56 1965 58
rect 1959 54 1961 56
rect 1963 54 1965 56
rect 1959 52 1965 54
rect 1963 49 1965 52
rect 1912 47 1914 49
rect 1916 47 1918 49
rect 1912 45 1918 47
rect 1896 27 1898 32
rect 1855 18 1857 22
rect 1876 18 1878 22
rect 1883 18 1885 22
rect 1943 27 1945 31
rect 1953 27 1955 31
rect 1927 18 1929 22
rect 1983 47 1985 60
rect 1993 56 1995 69
rect 1989 54 1995 56
rect 1989 52 1991 54
rect 1993 52 1995 54
rect 2003 59 2005 62
rect 2013 59 2015 62
rect 2033 59 2035 62
rect 2040 59 2042 62
rect 2051 59 2053 68
rect 2073 59 2075 68
rect 2111 76 2113 81
rect 2121 76 2123 81
rect 2131 79 2133 84
rect 2141 82 2143 86
rect 2206 84 2225 86
rect 2084 59 2086 62
rect 2091 59 2093 62
rect 2111 59 2113 62
rect 2121 59 2123 62
rect 2003 57 2009 59
rect 2003 55 2005 57
rect 2007 55 2009 57
rect 2003 53 2009 55
rect 2013 57 2035 59
rect 2013 55 2024 57
rect 2026 55 2031 57
rect 2033 55 2035 57
rect 2013 53 2035 55
rect 2039 57 2045 59
rect 2039 55 2041 57
rect 2043 55 2045 57
rect 2039 53 2045 55
rect 2049 57 2055 59
rect 2049 55 2051 57
rect 2053 55 2055 57
rect 2049 53 2055 55
rect 2071 57 2077 59
rect 2071 55 2073 57
rect 2075 55 2077 57
rect 2071 53 2077 55
rect 2081 57 2087 59
rect 2081 55 2083 57
rect 2085 55 2087 57
rect 2081 53 2087 55
rect 2091 57 2113 59
rect 2091 55 2093 57
rect 2095 55 2100 57
rect 2102 55 2113 57
rect 2091 53 2113 55
rect 2117 57 2123 59
rect 2117 55 2119 57
rect 2121 55 2123 57
rect 2117 53 2123 55
rect 2131 56 2133 69
rect 2141 66 2143 69
rect 2137 64 2143 66
rect 2137 62 2139 64
rect 2141 62 2143 64
rect 2162 68 2164 73
rect 2172 68 2174 73
rect 2182 71 2184 76
rect 2206 74 2208 84
rect 2216 76 2218 80
rect 2223 76 2225 84
rect 2274 84 2293 86
rect 2233 76 2235 81
rect 2240 76 2242 81
rect 2250 76 2252 81
rect 2137 60 2143 62
rect 2131 54 2137 56
rect 1989 50 1998 52
rect 2006 50 2008 53
rect 2013 50 2015 53
rect 2031 50 2033 53
rect 2041 50 2043 53
rect 2051 50 2053 53
rect 2073 50 2075 53
rect 2083 50 2085 53
rect 2093 50 2095 53
rect 2111 50 2113 53
rect 2118 50 2120 53
rect 2131 52 2133 54
rect 2135 52 2137 54
rect 2128 50 2137 52
rect 1996 47 1998 50
rect 1996 29 1998 34
rect 1963 18 1965 22
rect 1983 18 1985 22
rect 2006 20 2008 25
rect 2013 20 2015 25
rect 2128 47 2130 50
rect 2141 47 2143 60
rect 2162 52 2164 62
rect 2172 59 2174 62
rect 2182 59 2184 62
rect 2168 57 2174 59
rect 2168 55 2170 57
rect 2172 55 2174 57
rect 2168 53 2174 55
rect 2178 57 2184 59
rect 2178 55 2180 57
rect 2182 55 2184 57
rect 2178 53 2184 55
rect 2158 50 2164 52
rect 2158 48 2160 50
rect 2162 48 2164 50
rect 2128 29 2130 34
rect 2031 18 2033 22
rect 2041 18 2043 22
rect 2051 18 2053 22
rect 2073 18 2075 22
rect 2083 18 2085 22
rect 2093 18 2095 22
rect 2111 20 2113 25
rect 2118 20 2120 25
rect 2158 46 2164 48
rect 2162 43 2164 46
rect 2169 43 2171 53
rect 2182 50 2184 53
rect 2206 50 2208 68
rect 2216 59 2218 68
rect 2212 57 2218 59
rect 2212 55 2214 57
rect 2216 55 2218 57
rect 2212 53 2218 55
rect 2223 55 2225 68
rect 2233 65 2235 68
rect 2229 63 2235 65
rect 2229 61 2231 63
rect 2233 61 2235 63
rect 2229 59 2235 61
rect 2223 53 2235 55
rect 2240 54 2242 68
rect 2274 74 2276 84
rect 2284 76 2286 80
rect 2291 76 2293 84
rect 2301 76 2303 81
rect 2308 76 2310 81
rect 2318 76 2320 81
rect 2250 64 2252 67
rect 2247 62 2253 64
rect 2247 60 2249 62
rect 2251 60 2253 62
rect 2247 58 2253 60
rect 2206 39 2208 42
rect 2199 37 2208 39
rect 2216 38 2218 53
rect 2222 47 2228 49
rect 2222 45 2224 47
rect 2226 45 2228 47
rect 2222 43 2228 45
rect 2223 38 2225 43
rect 2233 38 2235 53
rect 2239 52 2245 54
rect 2239 50 2241 52
rect 2243 50 2245 52
rect 2239 48 2245 50
rect 2240 38 2242 48
rect 2250 40 2252 58
rect 2274 50 2276 68
rect 2284 59 2286 68
rect 2280 57 2286 59
rect 2280 55 2282 57
rect 2284 55 2286 57
rect 2280 53 2286 55
rect 2291 55 2293 68
rect 2301 65 2303 68
rect 2297 63 2303 65
rect 2297 61 2299 63
rect 2301 61 2303 63
rect 2297 59 2303 61
rect 2291 53 2303 55
rect 2308 54 2310 68
rect 2318 64 2320 67
rect 2315 62 2321 64
rect 2315 60 2317 62
rect 2319 60 2321 62
rect 2315 58 2321 60
rect 2199 35 2201 37
rect 2203 35 2205 37
rect 2199 33 2205 35
rect 2182 27 2184 32
rect 2141 18 2143 22
rect 2162 18 2164 22
rect 2169 18 2171 22
rect 2274 39 2276 42
rect 2267 37 2276 39
rect 2284 38 2286 53
rect 2290 47 2296 49
rect 2290 45 2292 47
rect 2294 45 2296 47
rect 2290 43 2296 45
rect 2291 38 2293 43
rect 2301 38 2303 53
rect 2307 52 2313 54
rect 2307 50 2309 52
rect 2311 50 2313 52
rect 2307 48 2313 50
rect 2308 38 2310 48
rect 2318 40 2320 58
rect 2267 35 2269 37
rect 2271 35 2273 37
rect 2267 33 2273 35
rect 2216 18 2218 22
rect 2223 18 2225 22
rect 2233 18 2235 22
rect 2240 18 2242 22
rect 2250 18 2252 22
rect 2284 18 2286 22
rect 2291 18 2293 22
rect 2301 18 2303 22
rect 2308 18 2310 22
rect 2318 18 2320 22
rect 15 3 17 8
rect 25 3 27 8
rect 95 10 97 14
rect 35 1 37 5
rect 55 3 57 8
rect 65 3 67 8
rect 15 -13 17 -10
rect 11 -15 17 -13
rect 11 -17 13 -15
rect 15 -17 17 -15
rect 11 -19 17 -17
rect 15 -32 17 -19
rect 25 -21 27 -10
rect 75 1 77 5
rect 55 -13 57 -10
rect 51 -15 57 -13
rect 51 -17 53 -15
rect 55 -17 57 -15
rect 35 -21 37 -17
rect 51 -19 57 -17
rect 21 -23 27 -21
rect 21 -25 23 -23
rect 25 -25 27 -23
rect 21 -27 27 -25
rect 31 -23 37 -21
rect 31 -25 33 -23
rect 35 -25 37 -23
rect 31 -27 37 -25
rect 22 -32 24 -27
rect 35 -32 37 -27
rect 55 -32 57 -19
rect 65 -21 67 -10
rect 118 7 120 12
rect 125 7 127 12
rect 143 10 145 14
rect 153 10 155 14
rect 163 10 165 14
rect 185 10 187 14
rect 195 10 197 14
rect 205 10 207 14
rect 108 -2 110 3
rect 75 -21 77 -17
rect 61 -23 67 -21
rect 61 -25 63 -23
rect 65 -25 67 -23
rect 61 -27 67 -25
rect 71 -23 77 -21
rect 71 -25 73 -23
rect 75 -25 77 -23
rect 71 -27 77 -25
rect 62 -32 64 -27
rect 75 -32 77 -27
rect 95 -28 97 -15
rect 108 -18 110 -15
rect 223 7 225 12
rect 230 7 232 12
rect 253 10 255 14
rect 274 10 276 14
rect 281 10 283 14
rect 240 -2 242 3
rect 362 10 364 14
rect 294 0 296 5
rect 322 3 324 8
rect 332 3 334 8
rect 274 -14 276 -11
rect 240 -18 242 -15
rect 101 -20 110 -18
rect 101 -22 103 -20
rect 105 -22 107 -20
rect 118 -21 120 -18
rect 125 -21 127 -18
rect 143 -21 145 -18
rect 153 -21 155 -18
rect 163 -21 165 -18
rect 185 -21 187 -18
rect 195 -21 197 -18
rect 205 -21 207 -18
rect 223 -21 225 -18
rect 230 -21 232 -18
rect 240 -20 249 -18
rect 101 -24 107 -22
rect 95 -30 101 -28
rect 95 -32 97 -30
rect 99 -32 101 -30
rect 15 -48 17 -43
rect 22 -48 24 -43
rect 35 -45 37 -41
rect 95 -34 101 -32
rect 95 -37 97 -34
rect 105 -37 107 -24
rect 115 -23 121 -21
rect 115 -25 117 -23
rect 119 -25 121 -23
rect 115 -27 121 -25
rect 125 -23 147 -21
rect 125 -25 136 -23
rect 138 -25 143 -23
rect 145 -25 147 -23
rect 125 -27 147 -25
rect 151 -23 157 -21
rect 151 -25 153 -23
rect 155 -25 157 -23
rect 151 -27 157 -25
rect 161 -23 167 -21
rect 161 -25 163 -23
rect 165 -25 167 -23
rect 161 -27 167 -25
rect 183 -23 189 -21
rect 183 -25 185 -23
rect 187 -25 189 -23
rect 183 -27 189 -25
rect 193 -23 199 -21
rect 193 -25 195 -23
rect 197 -25 199 -23
rect 193 -27 199 -25
rect 203 -23 225 -21
rect 203 -25 205 -23
rect 207 -25 212 -23
rect 214 -25 225 -23
rect 203 -27 225 -25
rect 229 -23 235 -21
rect 229 -25 231 -23
rect 233 -25 235 -23
rect 229 -27 235 -25
rect 115 -30 117 -27
rect 125 -30 127 -27
rect 145 -30 147 -27
rect 152 -30 154 -27
rect 55 -48 57 -43
rect 62 -48 64 -43
rect 75 -45 77 -41
rect 95 -54 97 -50
rect 105 -52 107 -47
rect 115 -49 117 -44
rect 125 -49 127 -44
rect 163 -36 165 -27
rect 185 -36 187 -27
rect 196 -30 198 -27
rect 203 -30 205 -27
rect 223 -30 225 -27
rect 233 -30 235 -27
rect 243 -22 245 -20
rect 247 -22 249 -20
rect 243 -24 249 -22
rect 243 -37 245 -24
rect 253 -28 255 -15
rect 270 -16 276 -14
rect 270 -18 272 -16
rect 274 -18 276 -16
rect 270 -20 276 -18
rect 249 -30 255 -28
rect 274 -30 276 -20
rect 281 -21 283 -11
rect 342 1 344 5
rect 322 -13 324 -10
rect 318 -15 324 -13
rect 318 -17 320 -15
rect 322 -17 324 -15
rect 294 -21 296 -18
rect 318 -19 324 -17
rect 280 -23 286 -21
rect 280 -25 282 -23
rect 284 -25 286 -23
rect 280 -27 286 -25
rect 290 -23 296 -21
rect 290 -25 292 -23
rect 294 -25 296 -23
rect 290 -27 296 -25
rect 284 -30 286 -27
rect 294 -30 296 -27
rect 249 -32 251 -30
rect 253 -32 255 -30
rect 249 -34 255 -32
rect 253 -37 255 -34
rect 223 -49 225 -44
rect 233 -49 235 -44
rect 145 -54 147 -50
rect 152 -54 154 -50
rect 163 -54 165 -50
rect 185 -54 187 -50
rect 196 -54 198 -50
rect 203 -54 205 -50
rect 243 -52 245 -47
rect 274 -41 276 -36
rect 284 -41 286 -36
rect 322 -32 324 -19
rect 332 -21 334 -10
rect 385 7 387 12
rect 392 7 394 12
rect 410 10 412 14
rect 420 10 422 14
rect 430 10 432 14
rect 452 10 454 14
rect 462 10 464 14
rect 472 10 474 14
rect 375 -2 377 3
rect 342 -21 344 -17
rect 328 -23 334 -21
rect 328 -25 330 -23
rect 332 -25 334 -23
rect 328 -27 334 -25
rect 338 -23 344 -21
rect 338 -25 340 -23
rect 342 -25 344 -23
rect 338 -27 344 -25
rect 329 -32 331 -27
rect 342 -32 344 -27
rect 362 -28 364 -15
rect 375 -18 377 -15
rect 490 7 492 12
rect 497 7 499 12
rect 520 10 522 14
rect 541 10 543 14
rect 548 10 550 14
rect 507 -2 509 3
rect 629 10 631 14
rect 561 0 563 5
rect 589 3 591 8
rect 599 3 601 8
rect 541 -14 543 -11
rect 507 -18 509 -15
rect 368 -20 377 -18
rect 368 -22 370 -20
rect 372 -22 374 -20
rect 385 -21 387 -18
rect 392 -21 394 -18
rect 410 -21 412 -18
rect 420 -21 422 -18
rect 430 -21 432 -18
rect 452 -21 454 -18
rect 462 -21 464 -18
rect 472 -21 474 -18
rect 490 -21 492 -18
rect 497 -21 499 -18
rect 507 -20 516 -18
rect 368 -24 374 -22
rect 362 -30 368 -28
rect 362 -32 364 -30
rect 366 -32 368 -30
rect 294 -44 296 -39
rect 362 -34 368 -32
rect 362 -37 364 -34
rect 372 -37 374 -24
rect 382 -23 388 -21
rect 382 -25 384 -23
rect 386 -25 388 -23
rect 382 -27 388 -25
rect 392 -23 414 -21
rect 392 -25 403 -23
rect 405 -25 410 -23
rect 412 -25 414 -23
rect 392 -27 414 -25
rect 418 -23 424 -21
rect 418 -25 420 -23
rect 422 -25 424 -23
rect 418 -27 424 -25
rect 428 -23 434 -21
rect 428 -25 430 -23
rect 432 -25 434 -23
rect 428 -27 434 -25
rect 450 -23 456 -21
rect 450 -25 452 -23
rect 454 -25 456 -23
rect 450 -27 456 -25
rect 460 -23 466 -21
rect 460 -25 462 -23
rect 464 -25 466 -23
rect 460 -27 466 -25
rect 470 -23 492 -21
rect 470 -25 472 -23
rect 474 -25 479 -23
rect 481 -25 492 -23
rect 470 -27 492 -25
rect 496 -23 502 -21
rect 496 -25 498 -23
rect 500 -25 502 -23
rect 496 -27 502 -25
rect 382 -30 384 -27
rect 392 -30 394 -27
rect 412 -30 414 -27
rect 419 -30 421 -27
rect 322 -48 324 -43
rect 329 -48 331 -43
rect 253 -54 255 -50
rect 342 -45 344 -41
rect 362 -54 364 -50
rect 372 -52 374 -47
rect 382 -49 384 -44
rect 392 -49 394 -44
rect 430 -36 432 -27
rect 452 -36 454 -27
rect 463 -30 465 -27
rect 470 -30 472 -27
rect 490 -30 492 -27
rect 500 -30 502 -27
rect 510 -22 512 -20
rect 514 -22 516 -20
rect 510 -24 516 -22
rect 510 -37 512 -24
rect 520 -28 522 -15
rect 537 -16 543 -14
rect 537 -18 539 -16
rect 541 -18 543 -16
rect 537 -20 543 -18
rect 516 -30 522 -28
rect 541 -30 543 -20
rect 548 -21 550 -11
rect 609 1 611 5
rect 589 -13 591 -10
rect 585 -15 591 -13
rect 585 -17 587 -15
rect 589 -17 591 -15
rect 561 -21 563 -18
rect 585 -19 591 -17
rect 547 -23 553 -21
rect 547 -25 549 -23
rect 551 -25 553 -23
rect 547 -27 553 -25
rect 557 -23 563 -21
rect 557 -25 559 -23
rect 561 -25 563 -23
rect 557 -27 563 -25
rect 551 -30 553 -27
rect 561 -30 563 -27
rect 516 -32 518 -30
rect 520 -32 522 -30
rect 516 -34 522 -32
rect 520 -37 522 -34
rect 490 -49 492 -44
rect 500 -49 502 -44
rect 412 -54 414 -50
rect 419 -54 421 -50
rect 430 -54 432 -50
rect 452 -54 454 -50
rect 463 -54 465 -50
rect 470 -54 472 -50
rect 510 -52 512 -47
rect 541 -41 543 -36
rect 551 -41 553 -36
rect 589 -32 591 -19
rect 599 -21 601 -10
rect 652 7 654 12
rect 659 7 661 12
rect 677 10 679 14
rect 687 10 689 14
rect 697 10 699 14
rect 719 10 721 14
rect 729 10 731 14
rect 739 10 741 14
rect 642 -2 644 3
rect 609 -21 611 -17
rect 595 -23 601 -21
rect 595 -25 597 -23
rect 599 -25 601 -23
rect 595 -27 601 -25
rect 605 -23 611 -21
rect 605 -25 607 -23
rect 609 -25 611 -23
rect 605 -27 611 -25
rect 596 -32 598 -27
rect 609 -32 611 -27
rect 629 -28 631 -15
rect 642 -18 644 -15
rect 757 7 759 12
rect 764 7 766 12
rect 787 10 789 14
rect 808 10 810 14
rect 815 10 817 14
rect 774 -2 776 3
rect 896 10 898 14
rect 828 0 830 5
rect 856 3 858 8
rect 866 3 868 8
rect 808 -14 810 -11
rect 774 -18 776 -15
rect 635 -20 644 -18
rect 635 -22 637 -20
rect 639 -22 641 -20
rect 652 -21 654 -18
rect 659 -21 661 -18
rect 677 -21 679 -18
rect 687 -21 689 -18
rect 697 -21 699 -18
rect 719 -21 721 -18
rect 729 -21 731 -18
rect 739 -21 741 -18
rect 757 -21 759 -18
rect 764 -21 766 -18
rect 774 -20 783 -18
rect 635 -24 641 -22
rect 629 -30 635 -28
rect 629 -32 631 -30
rect 633 -32 635 -30
rect 561 -44 563 -39
rect 629 -34 635 -32
rect 629 -37 631 -34
rect 639 -37 641 -24
rect 649 -23 655 -21
rect 649 -25 651 -23
rect 653 -25 655 -23
rect 649 -27 655 -25
rect 659 -23 681 -21
rect 659 -25 670 -23
rect 672 -25 677 -23
rect 679 -25 681 -23
rect 659 -27 681 -25
rect 685 -23 691 -21
rect 685 -25 687 -23
rect 689 -25 691 -23
rect 685 -27 691 -25
rect 695 -23 701 -21
rect 695 -25 697 -23
rect 699 -25 701 -23
rect 695 -27 701 -25
rect 717 -23 723 -21
rect 717 -25 719 -23
rect 721 -25 723 -23
rect 717 -27 723 -25
rect 727 -23 733 -21
rect 727 -25 729 -23
rect 731 -25 733 -23
rect 727 -27 733 -25
rect 737 -23 759 -21
rect 737 -25 739 -23
rect 741 -25 746 -23
rect 748 -25 759 -23
rect 737 -27 759 -25
rect 763 -23 769 -21
rect 763 -25 765 -23
rect 767 -25 769 -23
rect 763 -27 769 -25
rect 649 -30 651 -27
rect 659 -30 661 -27
rect 679 -30 681 -27
rect 686 -30 688 -27
rect 589 -48 591 -43
rect 596 -48 598 -43
rect 520 -54 522 -50
rect 609 -45 611 -41
rect 629 -54 631 -50
rect 639 -52 641 -47
rect 649 -49 651 -44
rect 659 -49 661 -44
rect 697 -36 699 -27
rect 719 -36 721 -27
rect 730 -30 732 -27
rect 737 -30 739 -27
rect 757 -30 759 -27
rect 767 -30 769 -27
rect 777 -22 779 -20
rect 781 -22 783 -20
rect 777 -24 783 -22
rect 777 -37 779 -24
rect 787 -28 789 -15
rect 804 -16 810 -14
rect 804 -18 806 -16
rect 808 -18 810 -16
rect 804 -20 810 -18
rect 783 -30 789 -28
rect 808 -30 810 -20
rect 815 -21 817 -11
rect 876 1 878 5
rect 856 -13 858 -10
rect 852 -15 858 -13
rect 852 -17 854 -15
rect 856 -17 858 -15
rect 828 -21 830 -18
rect 852 -19 858 -17
rect 814 -23 820 -21
rect 814 -25 816 -23
rect 818 -25 820 -23
rect 814 -27 820 -25
rect 824 -23 830 -21
rect 824 -25 826 -23
rect 828 -25 830 -23
rect 824 -27 830 -25
rect 818 -30 820 -27
rect 828 -30 830 -27
rect 783 -32 785 -30
rect 787 -32 789 -30
rect 783 -34 789 -32
rect 787 -37 789 -34
rect 757 -49 759 -44
rect 767 -49 769 -44
rect 679 -54 681 -50
rect 686 -54 688 -50
rect 697 -54 699 -50
rect 719 -54 721 -50
rect 730 -54 732 -50
rect 737 -54 739 -50
rect 777 -52 779 -47
rect 808 -41 810 -36
rect 818 -41 820 -36
rect 856 -32 858 -19
rect 866 -21 868 -10
rect 919 7 921 12
rect 926 7 928 12
rect 944 10 946 14
rect 954 10 956 14
rect 964 10 966 14
rect 986 10 988 14
rect 996 10 998 14
rect 1006 10 1008 14
rect 909 -2 911 3
rect 876 -21 878 -17
rect 862 -23 868 -21
rect 862 -25 864 -23
rect 866 -25 868 -23
rect 862 -27 868 -25
rect 872 -23 878 -21
rect 872 -25 874 -23
rect 876 -25 878 -23
rect 872 -27 878 -25
rect 863 -32 865 -27
rect 876 -32 878 -27
rect 896 -28 898 -15
rect 909 -18 911 -15
rect 1024 7 1026 12
rect 1031 7 1033 12
rect 1054 10 1056 14
rect 1075 10 1077 14
rect 1082 10 1084 14
rect 1041 -2 1043 3
rect 1163 10 1165 14
rect 1095 0 1097 5
rect 1123 3 1125 8
rect 1133 3 1135 8
rect 1075 -14 1077 -11
rect 1041 -18 1043 -15
rect 902 -20 911 -18
rect 902 -22 904 -20
rect 906 -22 908 -20
rect 919 -21 921 -18
rect 926 -21 928 -18
rect 944 -21 946 -18
rect 954 -21 956 -18
rect 964 -21 966 -18
rect 986 -21 988 -18
rect 996 -21 998 -18
rect 1006 -21 1008 -18
rect 1024 -21 1026 -18
rect 1031 -21 1033 -18
rect 1041 -20 1050 -18
rect 902 -24 908 -22
rect 896 -30 902 -28
rect 896 -32 898 -30
rect 900 -32 902 -30
rect 828 -44 830 -39
rect 896 -34 902 -32
rect 896 -37 898 -34
rect 906 -37 908 -24
rect 916 -23 922 -21
rect 916 -25 918 -23
rect 920 -25 922 -23
rect 916 -27 922 -25
rect 926 -23 948 -21
rect 926 -25 937 -23
rect 939 -25 944 -23
rect 946 -25 948 -23
rect 926 -27 948 -25
rect 952 -23 958 -21
rect 952 -25 954 -23
rect 956 -25 958 -23
rect 952 -27 958 -25
rect 962 -23 968 -21
rect 962 -25 964 -23
rect 966 -25 968 -23
rect 962 -27 968 -25
rect 984 -23 990 -21
rect 984 -25 986 -23
rect 988 -25 990 -23
rect 984 -27 990 -25
rect 994 -23 1000 -21
rect 994 -25 996 -23
rect 998 -25 1000 -23
rect 994 -27 1000 -25
rect 1004 -23 1026 -21
rect 1004 -25 1006 -23
rect 1008 -25 1013 -23
rect 1015 -25 1026 -23
rect 1004 -27 1026 -25
rect 1030 -23 1036 -21
rect 1030 -25 1032 -23
rect 1034 -25 1036 -23
rect 1030 -27 1036 -25
rect 916 -30 918 -27
rect 926 -30 928 -27
rect 946 -30 948 -27
rect 953 -30 955 -27
rect 856 -48 858 -43
rect 863 -48 865 -43
rect 787 -54 789 -50
rect 876 -45 878 -41
rect 896 -54 898 -50
rect 906 -52 908 -47
rect 916 -49 918 -44
rect 926 -49 928 -44
rect 964 -36 966 -27
rect 986 -36 988 -27
rect 997 -30 999 -27
rect 1004 -30 1006 -27
rect 1024 -30 1026 -27
rect 1034 -30 1036 -27
rect 1044 -22 1046 -20
rect 1048 -22 1050 -20
rect 1044 -24 1050 -22
rect 1044 -37 1046 -24
rect 1054 -28 1056 -15
rect 1071 -16 1077 -14
rect 1071 -18 1073 -16
rect 1075 -18 1077 -16
rect 1071 -20 1077 -18
rect 1050 -30 1056 -28
rect 1075 -30 1077 -20
rect 1082 -21 1084 -11
rect 1143 1 1145 5
rect 1123 -13 1125 -10
rect 1119 -15 1125 -13
rect 1119 -17 1121 -15
rect 1123 -17 1125 -15
rect 1095 -21 1097 -18
rect 1119 -19 1125 -17
rect 1081 -23 1087 -21
rect 1081 -25 1083 -23
rect 1085 -25 1087 -23
rect 1081 -27 1087 -25
rect 1091 -23 1097 -21
rect 1091 -25 1093 -23
rect 1095 -25 1097 -23
rect 1091 -27 1097 -25
rect 1085 -30 1087 -27
rect 1095 -30 1097 -27
rect 1050 -32 1052 -30
rect 1054 -32 1056 -30
rect 1050 -34 1056 -32
rect 1054 -37 1056 -34
rect 1024 -49 1026 -44
rect 1034 -49 1036 -44
rect 946 -54 948 -50
rect 953 -54 955 -50
rect 964 -54 966 -50
rect 986 -54 988 -50
rect 997 -54 999 -50
rect 1004 -54 1006 -50
rect 1044 -52 1046 -47
rect 1075 -41 1077 -36
rect 1085 -41 1087 -36
rect 1123 -32 1125 -19
rect 1133 -21 1135 -10
rect 1186 7 1188 12
rect 1193 7 1195 12
rect 1211 10 1213 14
rect 1221 10 1223 14
rect 1231 10 1233 14
rect 1253 10 1255 14
rect 1263 10 1265 14
rect 1273 10 1275 14
rect 1176 -2 1178 3
rect 1143 -21 1145 -17
rect 1129 -23 1135 -21
rect 1129 -25 1131 -23
rect 1133 -25 1135 -23
rect 1129 -27 1135 -25
rect 1139 -23 1145 -21
rect 1139 -25 1141 -23
rect 1143 -25 1145 -23
rect 1139 -27 1145 -25
rect 1130 -32 1132 -27
rect 1143 -32 1145 -27
rect 1163 -28 1165 -15
rect 1176 -18 1178 -15
rect 1291 7 1293 12
rect 1298 7 1300 12
rect 1321 10 1323 14
rect 1342 10 1344 14
rect 1349 10 1351 14
rect 1308 -2 1310 3
rect 1430 10 1432 14
rect 1362 0 1364 5
rect 1390 3 1392 8
rect 1400 3 1402 8
rect 1342 -14 1344 -11
rect 1308 -18 1310 -15
rect 1169 -20 1178 -18
rect 1169 -22 1171 -20
rect 1173 -22 1175 -20
rect 1186 -21 1188 -18
rect 1193 -21 1195 -18
rect 1211 -21 1213 -18
rect 1221 -21 1223 -18
rect 1231 -21 1233 -18
rect 1253 -21 1255 -18
rect 1263 -21 1265 -18
rect 1273 -21 1275 -18
rect 1291 -21 1293 -18
rect 1298 -21 1300 -18
rect 1308 -20 1317 -18
rect 1169 -24 1175 -22
rect 1163 -30 1169 -28
rect 1163 -32 1165 -30
rect 1167 -32 1169 -30
rect 1095 -44 1097 -39
rect 1163 -34 1169 -32
rect 1163 -37 1165 -34
rect 1173 -37 1175 -24
rect 1183 -23 1189 -21
rect 1183 -25 1185 -23
rect 1187 -25 1189 -23
rect 1183 -27 1189 -25
rect 1193 -23 1215 -21
rect 1193 -25 1204 -23
rect 1206 -25 1211 -23
rect 1213 -25 1215 -23
rect 1193 -27 1215 -25
rect 1219 -23 1225 -21
rect 1219 -25 1221 -23
rect 1223 -25 1225 -23
rect 1219 -27 1225 -25
rect 1229 -23 1235 -21
rect 1229 -25 1231 -23
rect 1233 -25 1235 -23
rect 1229 -27 1235 -25
rect 1251 -23 1257 -21
rect 1251 -25 1253 -23
rect 1255 -25 1257 -23
rect 1251 -27 1257 -25
rect 1261 -23 1267 -21
rect 1261 -25 1263 -23
rect 1265 -25 1267 -23
rect 1261 -27 1267 -25
rect 1271 -23 1293 -21
rect 1271 -25 1273 -23
rect 1275 -25 1280 -23
rect 1282 -25 1293 -23
rect 1271 -27 1293 -25
rect 1297 -23 1303 -21
rect 1297 -25 1299 -23
rect 1301 -25 1303 -23
rect 1297 -27 1303 -25
rect 1183 -30 1185 -27
rect 1193 -30 1195 -27
rect 1213 -30 1215 -27
rect 1220 -30 1222 -27
rect 1123 -48 1125 -43
rect 1130 -48 1132 -43
rect 1054 -54 1056 -50
rect 1143 -45 1145 -41
rect 1163 -54 1165 -50
rect 1173 -52 1175 -47
rect 1183 -49 1185 -44
rect 1193 -49 1195 -44
rect 1231 -36 1233 -27
rect 1253 -36 1255 -27
rect 1264 -30 1266 -27
rect 1271 -30 1273 -27
rect 1291 -30 1293 -27
rect 1301 -30 1303 -27
rect 1311 -22 1313 -20
rect 1315 -22 1317 -20
rect 1311 -24 1317 -22
rect 1311 -37 1313 -24
rect 1321 -28 1323 -15
rect 1338 -16 1344 -14
rect 1338 -18 1340 -16
rect 1342 -18 1344 -16
rect 1338 -20 1344 -18
rect 1317 -30 1323 -28
rect 1342 -30 1344 -20
rect 1349 -21 1351 -11
rect 1410 1 1412 5
rect 1390 -13 1392 -10
rect 1386 -15 1392 -13
rect 1386 -17 1388 -15
rect 1390 -17 1392 -15
rect 1362 -21 1364 -18
rect 1386 -19 1392 -17
rect 1348 -23 1354 -21
rect 1348 -25 1350 -23
rect 1352 -25 1354 -23
rect 1348 -27 1354 -25
rect 1358 -23 1364 -21
rect 1358 -25 1360 -23
rect 1362 -25 1364 -23
rect 1358 -27 1364 -25
rect 1352 -30 1354 -27
rect 1362 -30 1364 -27
rect 1317 -32 1319 -30
rect 1321 -32 1323 -30
rect 1317 -34 1323 -32
rect 1321 -37 1323 -34
rect 1291 -49 1293 -44
rect 1301 -49 1303 -44
rect 1213 -54 1215 -50
rect 1220 -54 1222 -50
rect 1231 -54 1233 -50
rect 1253 -54 1255 -50
rect 1264 -54 1266 -50
rect 1271 -54 1273 -50
rect 1311 -52 1313 -47
rect 1342 -41 1344 -36
rect 1352 -41 1354 -36
rect 1390 -32 1392 -19
rect 1400 -21 1402 -10
rect 1453 7 1455 12
rect 1460 7 1462 12
rect 1478 10 1480 14
rect 1488 10 1490 14
rect 1498 10 1500 14
rect 1520 10 1522 14
rect 1530 10 1532 14
rect 1540 10 1542 14
rect 1443 -2 1445 3
rect 1410 -21 1412 -17
rect 1396 -23 1402 -21
rect 1396 -25 1398 -23
rect 1400 -25 1402 -23
rect 1396 -27 1402 -25
rect 1406 -23 1412 -21
rect 1406 -25 1408 -23
rect 1410 -25 1412 -23
rect 1406 -27 1412 -25
rect 1397 -32 1399 -27
rect 1410 -32 1412 -27
rect 1430 -28 1432 -15
rect 1443 -18 1445 -15
rect 1558 7 1560 12
rect 1565 7 1567 12
rect 1588 10 1590 14
rect 1609 10 1611 14
rect 1616 10 1618 14
rect 1575 -2 1577 3
rect 1697 10 1699 14
rect 1629 0 1631 5
rect 1657 3 1659 8
rect 1667 3 1669 8
rect 1609 -14 1611 -11
rect 1575 -18 1577 -15
rect 1436 -20 1445 -18
rect 1436 -22 1438 -20
rect 1440 -22 1442 -20
rect 1453 -21 1455 -18
rect 1460 -21 1462 -18
rect 1478 -21 1480 -18
rect 1488 -21 1490 -18
rect 1498 -21 1500 -18
rect 1520 -21 1522 -18
rect 1530 -21 1532 -18
rect 1540 -21 1542 -18
rect 1558 -21 1560 -18
rect 1565 -21 1567 -18
rect 1575 -20 1584 -18
rect 1436 -24 1442 -22
rect 1430 -30 1436 -28
rect 1430 -32 1432 -30
rect 1434 -32 1436 -30
rect 1362 -44 1364 -39
rect 1430 -34 1436 -32
rect 1430 -37 1432 -34
rect 1440 -37 1442 -24
rect 1450 -23 1456 -21
rect 1450 -25 1452 -23
rect 1454 -25 1456 -23
rect 1450 -27 1456 -25
rect 1460 -23 1482 -21
rect 1460 -25 1471 -23
rect 1473 -25 1478 -23
rect 1480 -25 1482 -23
rect 1460 -27 1482 -25
rect 1486 -23 1492 -21
rect 1486 -25 1488 -23
rect 1490 -25 1492 -23
rect 1486 -27 1492 -25
rect 1496 -23 1502 -21
rect 1496 -25 1498 -23
rect 1500 -25 1502 -23
rect 1496 -27 1502 -25
rect 1518 -23 1524 -21
rect 1518 -25 1520 -23
rect 1522 -25 1524 -23
rect 1518 -27 1524 -25
rect 1528 -23 1534 -21
rect 1528 -25 1530 -23
rect 1532 -25 1534 -23
rect 1528 -27 1534 -25
rect 1538 -23 1560 -21
rect 1538 -25 1540 -23
rect 1542 -25 1547 -23
rect 1549 -25 1560 -23
rect 1538 -27 1560 -25
rect 1564 -23 1570 -21
rect 1564 -25 1566 -23
rect 1568 -25 1570 -23
rect 1564 -27 1570 -25
rect 1450 -30 1452 -27
rect 1460 -30 1462 -27
rect 1480 -30 1482 -27
rect 1487 -30 1489 -27
rect 1390 -48 1392 -43
rect 1397 -48 1399 -43
rect 1321 -54 1323 -50
rect 1410 -45 1412 -41
rect 1430 -54 1432 -50
rect 1440 -52 1442 -47
rect 1450 -49 1452 -44
rect 1460 -49 1462 -44
rect 1498 -36 1500 -27
rect 1520 -36 1522 -27
rect 1531 -30 1533 -27
rect 1538 -30 1540 -27
rect 1558 -30 1560 -27
rect 1568 -30 1570 -27
rect 1578 -22 1580 -20
rect 1582 -22 1584 -20
rect 1578 -24 1584 -22
rect 1578 -37 1580 -24
rect 1588 -28 1590 -15
rect 1605 -16 1611 -14
rect 1605 -18 1607 -16
rect 1609 -18 1611 -16
rect 1605 -20 1611 -18
rect 1584 -30 1590 -28
rect 1609 -30 1611 -20
rect 1616 -21 1618 -11
rect 1677 1 1679 5
rect 1657 -13 1659 -10
rect 1653 -15 1659 -13
rect 1653 -17 1655 -15
rect 1657 -17 1659 -15
rect 1629 -21 1631 -18
rect 1653 -19 1659 -17
rect 1615 -23 1621 -21
rect 1615 -25 1617 -23
rect 1619 -25 1621 -23
rect 1615 -27 1621 -25
rect 1625 -23 1631 -21
rect 1625 -25 1627 -23
rect 1629 -25 1631 -23
rect 1625 -27 1631 -25
rect 1619 -30 1621 -27
rect 1629 -30 1631 -27
rect 1584 -32 1586 -30
rect 1588 -32 1590 -30
rect 1584 -34 1590 -32
rect 1588 -37 1590 -34
rect 1558 -49 1560 -44
rect 1568 -49 1570 -44
rect 1480 -54 1482 -50
rect 1487 -54 1489 -50
rect 1498 -54 1500 -50
rect 1520 -54 1522 -50
rect 1531 -54 1533 -50
rect 1538 -54 1540 -50
rect 1578 -52 1580 -47
rect 1609 -41 1611 -36
rect 1619 -41 1621 -36
rect 1657 -32 1659 -19
rect 1667 -21 1669 -10
rect 1720 7 1722 12
rect 1727 7 1729 12
rect 1745 10 1747 14
rect 1755 10 1757 14
rect 1765 10 1767 14
rect 1787 10 1789 14
rect 1797 10 1799 14
rect 1807 10 1809 14
rect 1710 -2 1712 3
rect 1677 -21 1679 -17
rect 1663 -23 1669 -21
rect 1663 -25 1665 -23
rect 1667 -25 1669 -23
rect 1663 -27 1669 -25
rect 1673 -23 1679 -21
rect 1673 -25 1675 -23
rect 1677 -25 1679 -23
rect 1673 -27 1679 -25
rect 1664 -32 1666 -27
rect 1677 -32 1679 -27
rect 1697 -28 1699 -15
rect 1710 -18 1712 -15
rect 1825 7 1827 12
rect 1832 7 1834 12
rect 1855 10 1857 14
rect 1876 10 1878 14
rect 1883 10 1885 14
rect 1842 -2 1844 3
rect 1927 10 1929 14
rect 1896 0 1898 5
rect 1876 -14 1878 -11
rect 1842 -18 1844 -15
rect 1703 -20 1712 -18
rect 1703 -22 1705 -20
rect 1707 -22 1709 -20
rect 1720 -21 1722 -18
rect 1727 -21 1729 -18
rect 1745 -21 1747 -18
rect 1755 -21 1757 -18
rect 1765 -21 1767 -18
rect 1787 -21 1789 -18
rect 1797 -21 1799 -18
rect 1807 -21 1809 -18
rect 1825 -21 1827 -18
rect 1832 -21 1834 -18
rect 1842 -20 1851 -18
rect 1703 -24 1709 -22
rect 1697 -30 1703 -28
rect 1697 -32 1699 -30
rect 1701 -32 1703 -30
rect 1629 -44 1631 -39
rect 1697 -34 1703 -32
rect 1697 -37 1699 -34
rect 1707 -37 1709 -24
rect 1717 -23 1723 -21
rect 1717 -25 1719 -23
rect 1721 -25 1723 -23
rect 1717 -27 1723 -25
rect 1727 -23 1749 -21
rect 1727 -25 1738 -23
rect 1740 -25 1745 -23
rect 1747 -25 1749 -23
rect 1727 -27 1749 -25
rect 1753 -23 1759 -21
rect 1753 -25 1755 -23
rect 1757 -25 1759 -23
rect 1753 -27 1759 -25
rect 1763 -23 1769 -21
rect 1763 -25 1765 -23
rect 1767 -25 1769 -23
rect 1763 -27 1769 -25
rect 1785 -23 1791 -21
rect 1785 -25 1787 -23
rect 1789 -25 1791 -23
rect 1785 -27 1791 -25
rect 1795 -23 1801 -21
rect 1795 -25 1797 -23
rect 1799 -25 1801 -23
rect 1795 -27 1801 -25
rect 1805 -23 1827 -21
rect 1805 -25 1807 -23
rect 1809 -25 1814 -23
rect 1816 -25 1827 -23
rect 1805 -27 1827 -25
rect 1831 -23 1837 -21
rect 1831 -25 1833 -23
rect 1835 -25 1837 -23
rect 1831 -27 1837 -25
rect 1717 -30 1719 -27
rect 1727 -30 1729 -27
rect 1747 -30 1749 -27
rect 1754 -30 1756 -27
rect 1657 -48 1659 -43
rect 1664 -48 1666 -43
rect 1588 -54 1590 -50
rect 1677 -45 1679 -41
rect 1697 -54 1699 -50
rect 1707 -52 1709 -47
rect 1717 -49 1719 -44
rect 1727 -49 1729 -44
rect 1765 -36 1767 -27
rect 1787 -36 1789 -27
rect 1798 -30 1800 -27
rect 1805 -30 1807 -27
rect 1825 -30 1827 -27
rect 1835 -30 1837 -27
rect 1845 -22 1847 -20
rect 1849 -22 1851 -20
rect 1845 -24 1851 -22
rect 1845 -37 1847 -24
rect 1855 -28 1857 -15
rect 1872 -16 1878 -14
rect 1872 -18 1874 -16
rect 1876 -18 1878 -16
rect 1872 -20 1878 -18
rect 1851 -30 1857 -28
rect 1876 -30 1878 -20
rect 1883 -21 1885 -11
rect 1912 -15 1918 -13
rect 1912 -17 1914 -15
rect 1916 -17 1918 -15
rect 1963 10 1965 14
rect 1983 10 1985 14
rect 1943 1 1945 5
rect 1953 1 1955 5
rect 2006 7 2008 12
rect 2013 7 2015 12
rect 2031 10 2033 14
rect 2041 10 2043 14
rect 2051 10 2053 14
rect 2073 10 2075 14
rect 2083 10 2085 14
rect 2093 10 2095 14
rect 1996 -2 1998 3
rect 1896 -21 1898 -18
rect 1912 -19 1918 -17
rect 1882 -23 1888 -21
rect 1882 -25 1884 -23
rect 1886 -25 1888 -23
rect 1882 -27 1888 -25
rect 1892 -23 1898 -21
rect 1916 -20 1918 -19
rect 1927 -20 1929 -17
rect 1943 -20 1945 -17
rect 1916 -22 1929 -20
rect 1935 -22 1945 -20
rect 1953 -21 1955 -17
rect 1963 -20 1965 -17
rect 1892 -25 1894 -23
rect 1896 -25 1898 -23
rect 1892 -27 1898 -25
rect 1886 -30 1888 -27
rect 1896 -30 1898 -27
rect 1919 -30 1921 -22
rect 1935 -26 1937 -22
rect 1928 -28 1937 -26
rect 1949 -23 1955 -21
rect 1949 -25 1951 -23
rect 1953 -25 1955 -23
rect 1949 -27 1955 -25
rect 1959 -22 1965 -20
rect 1959 -24 1961 -22
rect 1963 -24 1965 -22
rect 1959 -26 1965 -24
rect 1928 -30 1930 -28
rect 1932 -30 1937 -28
rect 1851 -32 1853 -30
rect 1855 -32 1857 -30
rect 1851 -34 1857 -32
rect 1855 -37 1857 -34
rect 1825 -49 1827 -44
rect 1835 -49 1837 -44
rect 1747 -54 1749 -50
rect 1754 -54 1756 -50
rect 1765 -54 1767 -50
rect 1787 -54 1789 -50
rect 1798 -54 1800 -50
rect 1805 -54 1807 -50
rect 1845 -52 1847 -47
rect 1876 -41 1878 -36
rect 1886 -41 1888 -36
rect 1928 -32 1937 -30
rect 1953 -30 1955 -27
rect 1935 -35 1937 -32
rect 1945 -35 1947 -31
rect 1953 -32 1957 -30
rect 1955 -35 1957 -32
rect 1962 -35 1964 -26
rect 1983 -28 1985 -15
rect 1996 -18 1998 -15
rect 2111 7 2113 12
rect 2118 7 2120 12
rect 2141 10 2143 14
rect 2162 10 2164 14
rect 2169 10 2171 14
rect 2128 -2 2130 3
rect 2216 10 2218 14
rect 2223 10 2225 14
rect 2233 10 2235 14
rect 2240 10 2242 14
rect 2250 10 2252 14
rect 2284 10 2286 14
rect 2291 10 2293 14
rect 2301 10 2303 14
rect 2308 10 2310 14
rect 2318 10 2320 14
rect 2182 0 2184 5
rect 2162 -14 2164 -11
rect 2128 -18 2130 -15
rect 1989 -20 1998 -18
rect 1989 -22 1991 -20
rect 1993 -22 1995 -20
rect 2006 -21 2008 -18
rect 2013 -21 2015 -18
rect 2031 -21 2033 -18
rect 2041 -21 2043 -18
rect 2051 -21 2053 -18
rect 2073 -21 2075 -18
rect 2083 -21 2085 -18
rect 2093 -21 2095 -18
rect 2111 -21 2113 -18
rect 2118 -21 2120 -18
rect 2128 -20 2137 -18
rect 1989 -24 1995 -22
rect 1983 -30 1989 -28
rect 1983 -32 1985 -30
rect 1987 -32 1989 -30
rect 1983 -34 1989 -32
rect 1896 -44 1898 -39
rect 1919 -42 1921 -39
rect 1919 -44 1924 -42
rect 1855 -54 1857 -50
rect 1922 -52 1924 -44
rect 1935 -48 1937 -44
rect 1945 -52 1947 -44
rect 1983 -37 1985 -34
rect 1993 -37 1995 -24
rect 2003 -23 2009 -21
rect 2003 -25 2005 -23
rect 2007 -25 2009 -23
rect 2003 -27 2009 -25
rect 2013 -23 2035 -21
rect 2013 -25 2024 -23
rect 2026 -25 2031 -23
rect 2033 -25 2035 -23
rect 2013 -27 2035 -25
rect 2039 -23 2045 -21
rect 2039 -25 2041 -23
rect 2043 -25 2045 -23
rect 2039 -27 2045 -25
rect 2049 -23 2055 -21
rect 2049 -25 2051 -23
rect 2053 -25 2055 -23
rect 2049 -27 2055 -25
rect 2071 -23 2077 -21
rect 2071 -25 2073 -23
rect 2075 -25 2077 -23
rect 2071 -27 2077 -25
rect 2081 -23 2087 -21
rect 2081 -25 2083 -23
rect 2085 -25 2087 -23
rect 2081 -27 2087 -25
rect 2091 -23 2113 -21
rect 2091 -25 2093 -23
rect 2095 -25 2100 -23
rect 2102 -25 2113 -23
rect 2091 -27 2113 -25
rect 2117 -23 2123 -21
rect 2117 -25 2119 -23
rect 2121 -25 2123 -23
rect 2117 -27 2123 -25
rect 2003 -30 2005 -27
rect 2013 -30 2015 -27
rect 2033 -30 2035 -27
rect 2040 -30 2042 -27
rect 1955 -52 1957 -47
rect 1962 -52 1964 -47
rect 1922 -54 1947 -52
rect 1983 -54 1985 -50
rect 1993 -52 1995 -47
rect 2003 -49 2005 -44
rect 2013 -49 2015 -44
rect 2051 -36 2053 -27
rect 2073 -36 2075 -27
rect 2084 -30 2086 -27
rect 2091 -30 2093 -27
rect 2111 -30 2113 -27
rect 2121 -30 2123 -27
rect 2131 -22 2133 -20
rect 2135 -22 2137 -20
rect 2131 -24 2137 -22
rect 2131 -37 2133 -24
rect 2141 -28 2143 -15
rect 2158 -16 2164 -14
rect 2158 -18 2160 -16
rect 2162 -18 2164 -16
rect 2158 -20 2164 -18
rect 2137 -30 2143 -28
rect 2162 -30 2164 -20
rect 2169 -21 2171 -11
rect 2199 -3 2205 -1
rect 2199 -5 2201 -3
rect 2203 -5 2205 -3
rect 2199 -7 2208 -5
rect 2206 -10 2208 -7
rect 2182 -21 2184 -18
rect 2168 -23 2174 -21
rect 2168 -25 2170 -23
rect 2172 -25 2174 -23
rect 2168 -27 2174 -25
rect 2178 -23 2184 -21
rect 2178 -25 2180 -23
rect 2182 -25 2184 -23
rect 2178 -27 2184 -25
rect 2172 -30 2174 -27
rect 2182 -30 2184 -27
rect 2137 -32 2139 -30
rect 2141 -32 2143 -30
rect 2137 -34 2143 -32
rect 2141 -37 2143 -34
rect 2111 -49 2113 -44
rect 2121 -49 2123 -44
rect 2033 -54 2035 -50
rect 2040 -54 2042 -50
rect 2051 -54 2053 -50
rect 2073 -54 2075 -50
rect 2084 -54 2086 -50
rect 2091 -54 2093 -50
rect 2131 -52 2133 -47
rect 2162 -41 2164 -36
rect 2172 -41 2174 -36
rect 2206 -36 2208 -18
rect 2216 -21 2218 -6
rect 2223 -11 2225 -6
rect 2222 -13 2228 -11
rect 2222 -15 2224 -13
rect 2226 -15 2228 -13
rect 2222 -17 2228 -15
rect 2233 -21 2235 -6
rect 2240 -16 2242 -6
rect 2267 -3 2273 -1
rect 2267 -5 2269 -3
rect 2271 -5 2273 -3
rect 2267 -7 2276 -5
rect 2212 -23 2218 -21
rect 2212 -25 2214 -23
rect 2216 -25 2218 -23
rect 2212 -27 2218 -25
rect 2216 -36 2218 -27
rect 2223 -23 2235 -21
rect 2239 -18 2245 -16
rect 2239 -20 2241 -18
rect 2243 -20 2245 -18
rect 2239 -22 2245 -20
rect 2223 -36 2225 -23
rect 2229 -29 2235 -27
rect 2229 -31 2231 -29
rect 2233 -31 2235 -29
rect 2229 -33 2235 -31
rect 2233 -36 2235 -33
rect 2240 -36 2242 -22
rect 2250 -26 2252 -8
rect 2274 -10 2276 -7
rect 2247 -28 2253 -26
rect 2247 -30 2249 -28
rect 2251 -30 2253 -28
rect 2247 -32 2253 -30
rect 2250 -35 2252 -32
rect 2182 -44 2184 -39
rect 2141 -54 2143 -50
rect 2206 -52 2208 -42
rect 2274 -36 2276 -18
rect 2284 -21 2286 -6
rect 2291 -11 2293 -6
rect 2290 -13 2296 -11
rect 2290 -15 2292 -13
rect 2294 -15 2296 -13
rect 2290 -17 2296 -15
rect 2301 -21 2303 -6
rect 2308 -16 2310 -6
rect 2280 -23 2286 -21
rect 2280 -25 2282 -23
rect 2284 -25 2286 -23
rect 2280 -27 2286 -25
rect 2284 -36 2286 -27
rect 2291 -23 2303 -21
rect 2307 -18 2313 -16
rect 2307 -20 2309 -18
rect 2311 -20 2313 -18
rect 2307 -22 2313 -20
rect 2291 -36 2293 -23
rect 2297 -29 2303 -27
rect 2297 -31 2299 -29
rect 2301 -31 2303 -29
rect 2297 -33 2303 -31
rect 2301 -36 2303 -33
rect 2308 -36 2310 -22
rect 2318 -26 2320 -8
rect 2315 -28 2321 -26
rect 2315 -30 2317 -28
rect 2319 -30 2321 -28
rect 2315 -32 2321 -30
rect 2318 -35 2320 -32
rect 2216 -48 2218 -44
rect 2223 -52 2225 -44
rect 2233 -49 2235 -44
rect 2240 -49 2242 -44
rect 2250 -49 2252 -44
rect 2206 -54 2225 -52
rect 2274 -52 2276 -42
rect 2284 -48 2286 -44
rect 2291 -52 2293 -44
rect 2301 -49 2303 -44
rect 2308 -49 2310 -44
rect 2318 -49 2320 -44
rect 2274 -54 2293 -52
rect 15 -69 17 -64
rect 22 -69 24 -64
rect 35 -71 37 -67
rect 55 -69 57 -64
rect 62 -69 64 -64
rect 95 -62 97 -58
rect 75 -71 77 -67
rect 105 -65 107 -60
rect 145 -62 147 -58
rect 152 -62 154 -58
rect 163 -62 165 -58
rect 185 -62 187 -58
rect 196 -62 198 -58
rect 203 -62 205 -58
rect 115 -68 117 -63
rect 125 -68 127 -63
rect 95 -78 97 -75
rect 95 -80 101 -78
rect 15 -93 17 -80
rect 22 -85 24 -80
rect 35 -85 37 -80
rect 21 -87 27 -85
rect 21 -89 23 -87
rect 25 -89 27 -87
rect 21 -91 27 -89
rect 31 -87 37 -85
rect 31 -89 33 -87
rect 35 -89 37 -87
rect 31 -91 37 -89
rect 11 -95 17 -93
rect 11 -97 13 -95
rect 15 -97 17 -95
rect 11 -99 17 -97
rect 15 -102 17 -99
rect 25 -102 27 -91
rect 35 -95 37 -91
rect 55 -93 57 -80
rect 62 -85 64 -80
rect 75 -85 77 -80
rect 61 -87 67 -85
rect 61 -89 63 -87
rect 65 -89 67 -87
rect 61 -91 67 -89
rect 71 -87 77 -85
rect 71 -89 73 -87
rect 75 -89 77 -87
rect 71 -91 77 -89
rect 51 -95 57 -93
rect 51 -97 53 -95
rect 55 -97 57 -95
rect 51 -99 57 -97
rect 55 -102 57 -99
rect 65 -102 67 -91
rect 75 -95 77 -91
rect 95 -82 97 -80
rect 99 -82 101 -80
rect 95 -84 101 -82
rect 15 -120 17 -115
rect 25 -120 27 -115
rect 35 -117 37 -113
rect 95 -97 97 -84
rect 105 -88 107 -75
rect 101 -90 107 -88
rect 101 -92 103 -90
rect 105 -92 107 -90
rect 115 -85 117 -82
rect 125 -85 127 -82
rect 145 -85 147 -82
rect 152 -85 154 -82
rect 163 -85 165 -76
rect 185 -85 187 -76
rect 223 -68 225 -63
rect 233 -68 235 -63
rect 243 -65 245 -60
rect 253 -62 255 -58
rect 196 -85 198 -82
rect 203 -85 205 -82
rect 223 -85 225 -82
rect 233 -85 235 -82
rect 115 -87 121 -85
rect 115 -89 117 -87
rect 119 -89 121 -87
rect 115 -91 121 -89
rect 125 -87 147 -85
rect 125 -89 136 -87
rect 138 -89 143 -87
rect 145 -89 147 -87
rect 125 -91 147 -89
rect 151 -87 157 -85
rect 151 -89 153 -87
rect 155 -89 157 -87
rect 151 -91 157 -89
rect 161 -87 167 -85
rect 161 -89 163 -87
rect 165 -89 167 -87
rect 161 -91 167 -89
rect 183 -87 189 -85
rect 183 -89 185 -87
rect 187 -89 189 -87
rect 183 -91 189 -89
rect 193 -87 199 -85
rect 193 -89 195 -87
rect 197 -89 199 -87
rect 193 -91 199 -89
rect 203 -87 225 -85
rect 203 -89 205 -87
rect 207 -89 212 -87
rect 214 -89 225 -87
rect 203 -91 225 -89
rect 229 -87 235 -85
rect 229 -89 231 -87
rect 233 -89 235 -87
rect 229 -91 235 -89
rect 243 -88 245 -75
rect 253 -78 255 -75
rect 249 -80 255 -78
rect 249 -82 251 -80
rect 253 -82 255 -80
rect 274 -76 276 -71
rect 284 -76 286 -71
rect 294 -73 296 -68
rect 322 -69 324 -64
rect 329 -69 331 -64
rect 362 -62 364 -58
rect 342 -71 344 -67
rect 372 -65 374 -60
rect 412 -62 414 -58
rect 419 -62 421 -58
rect 430 -62 432 -58
rect 452 -62 454 -58
rect 463 -62 465 -58
rect 470 -62 472 -58
rect 382 -68 384 -63
rect 392 -68 394 -63
rect 362 -78 364 -75
rect 362 -80 368 -78
rect 249 -84 255 -82
rect 243 -90 249 -88
rect 101 -94 110 -92
rect 118 -94 120 -91
rect 125 -94 127 -91
rect 143 -94 145 -91
rect 153 -94 155 -91
rect 163 -94 165 -91
rect 185 -94 187 -91
rect 195 -94 197 -91
rect 205 -94 207 -91
rect 223 -94 225 -91
rect 230 -94 232 -91
rect 243 -92 245 -90
rect 247 -92 249 -90
rect 240 -94 249 -92
rect 108 -97 110 -94
rect 55 -120 57 -115
rect 65 -120 67 -115
rect 75 -117 77 -113
rect 108 -115 110 -110
rect 95 -126 97 -122
rect 118 -124 120 -119
rect 125 -124 127 -119
rect 240 -97 242 -94
rect 253 -97 255 -84
rect 274 -92 276 -82
rect 284 -85 286 -82
rect 294 -85 296 -82
rect 280 -87 286 -85
rect 280 -89 282 -87
rect 284 -89 286 -87
rect 280 -91 286 -89
rect 290 -87 296 -85
rect 290 -89 292 -87
rect 294 -89 296 -87
rect 290 -91 296 -89
rect 270 -94 276 -92
rect 270 -96 272 -94
rect 274 -96 276 -94
rect 240 -115 242 -110
rect 143 -126 145 -122
rect 153 -126 155 -122
rect 163 -126 165 -122
rect 185 -126 187 -122
rect 195 -126 197 -122
rect 205 -126 207 -122
rect 223 -124 225 -119
rect 230 -124 232 -119
rect 270 -98 276 -96
rect 274 -101 276 -98
rect 281 -101 283 -91
rect 294 -94 296 -91
rect 322 -93 324 -80
rect 329 -85 331 -80
rect 342 -85 344 -80
rect 328 -87 334 -85
rect 328 -89 330 -87
rect 332 -89 334 -87
rect 328 -91 334 -89
rect 338 -87 344 -85
rect 338 -89 340 -87
rect 342 -89 344 -87
rect 338 -91 344 -89
rect 318 -95 324 -93
rect 318 -97 320 -95
rect 322 -97 324 -95
rect 318 -99 324 -97
rect 322 -102 324 -99
rect 332 -102 334 -91
rect 342 -95 344 -91
rect 362 -82 364 -80
rect 366 -82 368 -80
rect 362 -84 368 -82
rect 294 -117 296 -112
rect 362 -97 364 -84
rect 372 -88 374 -75
rect 368 -90 374 -88
rect 368 -92 370 -90
rect 372 -92 374 -90
rect 382 -85 384 -82
rect 392 -85 394 -82
rect 412 -85 414 -82
rect 419 -85 421 -82
rect 430 -85 432 -76
rect 452 -85 454 -76
rect 490 -68 492 -63
rect 500 -68 502 -63
rect 510 -65 512 -60
rect 520 -62 522 -58
rect 463 -85 465 -82
rect 470 -85 472 -82
rect 490 -85 492 -82
rect 500 -85 502 -82
rect 382 -87 388 -85
rect 382 -89 384 -87
rect 386 -89 388 -87
rect 382 -91 388 -89
rect 392 -87 414 -85
rect 392 -89 403 -87
rect 405 -89 410 -87
rect 412 -89 414 -87
rect 392 -91 414 -89
rect 418 -87 424 -85
rect 418 -89 420 -87
rect 422 -89 424 -87
rect 418 -91 424 -89
rect 428 -87 434 -85
rect 428 -89 430 -87
rect 432 -89 434 -87
rect 428 -91 434 -89
rect 450 -87 456 -85
rect 450 -89 452 -87
rect 454 -89 456 -87
rect 450 -91 456 -89
rect 460 -87 466 -85
rect 460 -89 462 -87
rect 464 -89 466 -87
rect 460 -91 466 -89
rect 470 -87 492 -85
rect 470 -89 472 -87
rect 474 -89 479 -87
rect 481 -89 492 -87
rect 470 -91 492 -89
rect 496 -87 502 -85
rect 496 -89 498 -87
rect 500 -89 502 -87
rect 496 -91 502 -89
rect 510 -88 512 -75
rect 520 -78 522 -75
rect 516 -80 522 -78
rect 516 -82 518 -80
rect 520 -82 522 -80
rect 541 -76 543 -71
rect 551 -76 553 -71
rect 561 -73 563 -68
rect 589 -69 591 -64
rect 596 -69 598 -64
rect 629 -62 631 -58
rect 609 -71 611 -67
rect 639 -65 641 -60
rect 679 -62 681 -58
rect 686 -62 688 -58
rect 697 -62 699 -58
rect 719 -62 721 -58
rect 730 -62 732 -58
rect 737 -62 739 -58
rect 649 -68 651 -63
rect 659 -68 661 -63
rect 629 -78 631 -75
rect 629 -80 635 -78
rect 516 -84 522 -82
rect 510 -90 516 -88
rect 368 -94 377 -92
rect 385 -94 387 -91
rect 392 -94 394 -91
rect 410 -94 412 -91
rect 420 -94 422 -91
rect 430 -94 432 -91
rect 452 -94 454 -91
rect 462 -94 464 -91
rect 472 -94 474 -91
rect 490 -94 492 -91
rect 497 -94 499 -91
rect 510 -92 512 -90
rect 514 -92 516 -90
rect 507 -94 516 -92
rect 375 -97 377 -94
rect 322 -120 324 -115
rect 332 -120 334 -115
rect 342 -117 344 -113
rect 253 -126 255 -122
rect 274 -126 276 -122
rect 281 -126 283 -122
rect 375 -115 377 -110
rect 362 -126 364 -122
rect 385 -124 387 -119
rect 392 -124 394 -119
rect 507 -97 509 -94
rect 520 -97 522 -84
rect 541 -92 543 -82
rect 551 -85 553 -82
rect 561 -85 563 -82
rect 547 -87 553 -85
rect 547 -89 549 -87
rect 551 -89 553 -87
rect 547 -91 553 -89
rect 557 -87 563 -85
rect 557 -89 559 -87
rect 561 -89 563 -87
rect 557 -91 563 -89
rect 537 -94 543 -92
rect 537 -96 539 -94
rect 541 -96 543 -94
rect 507 -115 509 -110
rect 410 -126 412 -122
rect 420 -126 422 -122
rect 430 -126 432 -122
rect 452 -126 454 -122
rect 462 -126 464 -122
rect 472 -126 474 -122
rect 490 -124 492 -119
rect 497 -124 499 -119
rect 537 -98 543 -96
rect 541 -101 543 -98
rect 548 -101 550 -91
rect 561 -94 563 -91
rect 589 -93 591 -80
rect 596 -85 598 -80
rect 609 -85 611 -80
rect 595 -87 601 -85
rect 595 -89 597 -87
rect 599 -89 601 -87
rect 595 -91 601 -89
rect 605 -87 611 -85
rect 605 -89 607 -87
rect 609 -89 611 -87
rect 605 -91 611 -89
rect 585 -95 591 -93
rect 585 -97 587 -95
rect 589 -97 591 -95
rect 585 -99 591 -97
rect 589 -102 591 -99
rect 599 -102 601 -91
rect 609 -95 611 -91
rect 629 -82 631 -80
rect 633 -82 635 -80
rect 629 -84 635 -82
rect 561 -117 563 -112
rect 629 -97 631 -84
rect 639 -88 641 -75
rect 635 -90 641 -88
rect 635 -92 637 -90
rect 639 -92 641 -90
rect 649 -85 651 -82
rect 659 -85 661 -82
rect 679 -85 681 -82
rect 686 -85 688 -82
rect 697 -85 699 -76
rect 719 -85 721 -76
rect 757 -68 759 -63
rect 767 -68 769 -63
rect 777 -65 779 -60
rect 787 -62 789 -58
rect 730 -85 732 -82
rect 737 -85 739 -82
rect 757 -85 759 -82
rect 767 -85 769 -82
rect 649 -87 655 -85
rect 649 -89 651 -87
rect 653 -89 655 -87
rect 649 -91 655 -89
rect 659 -87 681 -85
rect 659 -89 670 -87
rect 672 -89 677 -87
rect 679 -89 681 -87
rect 659 -91 681 -89
rect 685 -87 691 -85
rect 685 -89 687 -87
rect 689 -89 691 -87
rect 685 -91 691 -89
rect 695 -87 701 -85
rect 695 -89 697 -87
rect 699 -89 701 -87
rect 695 -91 701 -89
rect 717 -87 723 -85
rect 717 -89 719 -87
rect 721 -89 723 -87
rect 717 -91 723 -89
rect 727 -87 733 -85
rect 727 -89 729 -87
rect 731 -89 733 -87
rect 727 -91 733 -89
rect 737 -87 759 -85
rect 737 -89 739 -87
rect 741 -89 746 -87
rect 748 -89 759 -87
rect 737 -91 759 -89
rect 763 -87 769 -85
rect 763 -89 765 -87
rect 767 -89 769 -87
rect 763 -91 769 -89
rect 777 -88 779 -75
rect 787 -78 789 -75
rect 783 -80 789 -78
rect 783 -82 785 -80
rect 787 -82 789 -80
rect 808 -76 810 -71
rect 818 -76 820 -71
rect 828 -73 830 -68
rect 856 -69 858 -64
rect 863 -69 865 -64
rect 896 -62 898 -58
rect 876 -71 878 -67
rect 906 -65 908 -60
rect 946 -62 948 -58
rect 953 -62 955 -58
rect 964 -62 966 -58
rect 986 -62 988 -58
rect 997 -62 999 -58
rect 1004 -62 1006 -58
rect 916 -68 918 -63
rect 926 -68 928 -63
rect 896 -78 898 -75
rect 896 -80 902 -78
rect 783 -84 789 -82
rect 777 -90 783 -88
rect 635 -94 644 -92
rect 652 -94 654 -91
rect 659 -94 661 -91
rect 677 -94 679 -91
rect 687 -94 689 -91
rect 697 -94 699 -91
rect 719 -94 721 -91
rect 729 -94 731 -91
rect 739 -94 741 -91
rect 757 -94 759 -91
rect 764 -94 766 -91
rect 777 -92 779 -90
rect 781 -92 783 -90
rect 774 -94 783 -92
rect 642 -97 644 -94
rect 589 -120 591 -115
rect 599 -120 601 -115
rect 609 -117 611 -113
rect 520 -126 522 -122
rect 541 -126 543 -122
rect 548 -126 550 -122
rect 642 -115 644 -110
rect 629 -126 631 -122
rect 652 -124 654 -119
rect 659 -124 661 -119
rect 774 -97 776 -94
rect 787 -97 789 -84
rect 808 -92 810 -82
rect 818 -85 820 -82
rect 828 -85 830 -82
rect 814 -87 820 -85
rect 814 -89 816 -87
rect 818 -89 820 -87
rect 814 -91 820 -89
rect 824 -87 830 -85
rect 824 -89 826 -87
rect 828 -89 830 -87
rect 824 -91 830 -89
rect 804 -94 810 -92
rect 804 -96 806 -94
rect 808 -96 810 -94
rect 774 -115 776 -110
rect 677 -126 679 -122
rect 687 -126 689 -122
rect 697 -126 699 -122
rect 719 -126 721 -122
rect 729 -126 731 -122
rect 739 -126 741 -122
rect 757 -124 759 -119
rect 764 -124 766 -119
rect 804 -98 810 -96
rect 808 -101 810 -98
rect 815 -101 817 -91
rect 828 -94 830 -91
rect 856 -93 858 -80
rect 863 -85 865 -80
rect 876 -85 878 -80
rect 862 -87 868 -85
rect 862 -89 864 -87
rect 866 -89 868 -87
rect 862 -91 868 -89
rect 872 -87 878 -85
rect 872 -89 874 -87
rect 876 -89 878 -87
rect 872 -91 878 -89
rect 852 -95 858 -93
rect 852 -97 854 -95
rect 856 -97 858 -95
rect 852 -99 858 -97
rect 856 -102 858 -99
rect 866 -102 868 -91
rect 876 -95 878 -91
rect 896 -82 898 -80
rect 900 -82 902 -80
rect 896 -84 902 -82
rect 828 -117 830 -112
rect 896 -97 898 -84
rect 906 -88 908 -75
rect 902 -90 908 -88
rect 902 -92 904 -90
rect 906 -92 908 -90
rect 916 -85 918 -82
rect 926 -85 928 -82
rect 946 -85 948 -82
rect 953 -85 955 -82
rect 964 -85 966 -76
rect 986 -85 988 -76
rect 1024 -68 1026 -63
rect 1034 -68 1036 -63
rect 1044 -65 1046 -60
rect 1054 -62 1056 -58
rect 997 -85 999 -82
rect 1004 -85 1006 -82
rect 1024 -85 1026 -82
rect 1034 -85 1036 -82
rect 916 -87 922 -85
rect 916 -89 918 -87
rect 920 -89 922 -87
rect 916 -91 922 -89
rect 926 -87 948 -85
rect 926 -89 937 -87
rect 939 -89 944 -87
rect 946 -89 948 -87
rect 926 -91 948 -89
rect 952 -87 958 -85
rect 952 -89 954 -87
rect 956 -89 958 -87
rect 952 -91 958 -89
rect 962 -87 968 -85
rect 962 -89 964 -87
rect 966 -89 968 -87
rect 962 -91 968 -89
rect 984 -87 990 -85
rect 984 -89 986 -87
rect 988 -89 990 -87
rect 984 -91 990 -89
rect 994 -87 1000 -85
rect 994 -89 996 -87
rect 998 -89 1000 -87
rect 994 -91 1000 -89
rect 1004 -87 1026 -85
rect 1004 -89 1006 -87
rect 1008 -89 1013 -87
rect 1015 -89 1026 -87
rect 1004 -91 1026 -89
rect 1030 -87 1036 -85
rect 1030 -89 1032 -87
rect 1034 -89 1036 -87
rect 1030 -91 1036 -89
rect 1044 -88 1046 -75
rect 1054 -78 1056 -75
rect 1050 -80 1056 -78
rect 1050 -82 1052 -80
rect 1054 -82 1056 -80
rect 1075 -76 1077 -71
rect 1085 -76 1087 -71
rect 1095 -73 1097 -68
rect 1123 -69 1125 -64
rect 1130 -69 1132 -64
rect 1163 -62 1165 -58
rect 1143 -71 1145 -67
rect 1173 -65 1175 -60
rect 1213 -62 1215 -58
rect 1220 -62 1222 -58
rect 1231 -62 1233 -58
rect 1253 -62 1255 -58
rect 1264 -62 1266 -58
rect 1271 -62 1273 -58
rect 1183 -68 1185 -63
rect 1193 -68 1195 -63
rect 1163 -78 1165 -75
rect 1163 -80 1169 -78
rect 1050 -84 1056 -82
rect 1044 -90 1050 -88
rect 902 -94 911 -92
rect 919 -94 921 -91
rect 926 -94 928 -91
rect 944 -94 946 -91
rect 954 -94 956 -91
rect 964 -94 966 -91
rect 986 -94 988 -91
rect 996 -94 998 -91
rect 1006 -94 1008 -91
rect 1024 -94 1026 -91
rect 1031 -94 1033 -91
rect 1044 -92 1046 -90
rect 1048 -92 1050 -90
rect 1041 -94 1050 -92
rect 909 -97 911 -94
rect 856 -120 858 -115
rect 866 -120 868 -115
rect 876 -117 878 -113
rect 787 -126 789 -122
rect 808 -126 810 -122
rect 815 -126 817 -122
rect 909 -115 911 -110
rect 896 -126 898 -122
rect 919 -124 921 -119
rect 926 -124 928 -119
rect 1041 -97 1043 -94
rect 1054 -97 1056 -84
rect 1075 -92 1077 -82
rect 1085 -85 1087 -82
rect 1095 -85 1097 -82
rect 1081 -87 1087 -85
rect 1081 -89 1083 -87
rect 1085 -89 1087 -87
rect 1081 -91 1087 -89
rect 1091 -87 1097 -85
rect 1091 -89 1093 -87
rect 1095 -89 1097 -87
rect 1091 -91 1097 -89
rect 1071 -94 1077 -92
rect 1071 -96 1073 -94
rect 1075 -96 1077 -94
rect 1041 -115 1043 -110
rect 944 -126 946 -122
rect 954 -126 956 -122
rect 964 -126 966 -122
rect 986 -126 988 -122
rect 996 -126 998 -122
rect 1006 -126 1008 -122
rect 1024 -124 1026 -119
rect 1031 -124 1033 -119
rect 1071 -98 1077 -96
rect 1075 -101 1077 -98
rect 1082 -101 1084 -91
rect 1095 -94 1097 -91
rect 1123 -93 1125 -80
rect 1130 -85 1132 -80
rect 1143 -85 1145 -80
rect 1129 -87 1135 -85
rect 1129 -89 1131 -87
rect 1133 -89 1135 -87
rect 1129 -91 1135 -89
rect 1139 -87 1145 -85
rect 1139 -89 1141 -87
rect 1143 -89 1145 -87
rect 1139 -91 1145 -89
rect 1119 -95 1125 -93
rect 1119 -97 1121 -95
rect 1123 -97 1125 -95
rect 1119 -99 1125 -97
rect 1123 -102 1125 -99
rect 1133 -102 1135 -91
rect 1143 -95 1145 -91
rect 1163 -82 1165 -80
rect 1167 -82 1169 -80
rect 1163 -84 1169 -82
rect 1095 -117 1097 -112
rect 1163 -97 1165 -84
rect 1173 -88 1175 -75
rect 1169 -90 1175 -88
rect 1169 -92 1171 -90
rect 1173 -92 1175 -90
rect 1183 -85 1185 -82
rect 1193 -85 1195 -82
rect 1213 -85 1215 -82
rect 1220 -85 1222 -82
rect 1231 -85 1233 -76
rect 1253 -85 1255 -76
rect 1291 -68 1293 -63
rect 1301 -68 1303 -63
rect 1311 -65 1313 -60
rect 1321 -62 1323 -58
rect 1264 -85 1266 -82
rect 1271 -85 1273 -82
rect 1291 -85 1293 -82
rect 1301 -85 1303 -82
rect 1183 -87 1189 -85
rect 1183 -89 1185 -87
rect 1187 -89 1189 -87
rect 1183 -91 1189 -89
rect 1193 -87 1215 -85
rect 1193 -89 1204 -87
rect 1206 -89 1211 -87
rect 1213 -89 1215 -87
rect 1193 -91 1215 -89
rect 1219 -87 1225 -85
rect 1219 -89 1221 -87
rect 1223 -89 1225 -87
rect 1219 -91 1225 -89
rect 1229 -87 1235 -85
rect 1229 -89 1231 -87
rect 1233 -89 1235 -87
rect 1229 -91 1235 -89
rect 1251 -87 1257 -85
rect 1251 -89 1253 -87
rect 1255 -89 1257 -87
rect 1251 -91 1257 -89
rect 1261 -87 1267 -85
rect 1261 -89 1263 -87
rect 1265 -89 1267 -87
rect 1261 -91 1267 -89
rect 1271 -87 1293 -85
rect 1271 -89 1273 -87
rect 1275 -89 1280 -87
rect 1282 -89 1293 -87
rect 1271 -91 1293 -89
rect 1297 -87 1303 -85
rect 1297 -89 1299 -87
rect 1301 -89 1303 -87
rect 1297 -91 1303 -89
rect 1311 -88 1313 -75
rect 1321 -78 1323 -75
rect 1317 -80 1323 -78
rect 1317 -82 1319 -80
rect 1321 -82 1323 -80
rect 1342 -76 1344 -71
rect 1352 -76 1354 -71
rect 1362 -73 1364 -68
rect 1390 -69 1392 -64
rect 1397 -69 1399 -64
rect 1430 -62 1432 -58
rect 1410 -71 1412 -67
rect 1440 -65 1442 -60
rect 1480 -62 1482 -58
rect 1487 -62 1489 -58
rect 1498 -62 1500 -58
rect 1520 -62 1522 -58
rect 1531 -62 1533 -58
rect 1538 -62 1540 -58
rect 1450 -68 1452 -63
rect 1460 -68 1462 -63
rect 1430 -78 1432 -75
rect 1430 -80 1436 -78
rect 1317 -84 1323 -82
rect 1311 -90 1317 -88
rect 1169 -94 1178 -92
rect 1186 -94 1188 -91
rect 1193 -94 1195 -91
rect 1211 -94 1213 -91
rect 1221 -94 1223 -91
rect 1231 -94 1233 -91
rect 1253 -94 1255 -91
rect 1263 -94 1265 -91
rect 1273 -94 1275 -91
rect 1291 -94 1293 -91
rect 1298 -94 1300 -91
rect 1311 -92 1313 -90
rect 1315 -92 1317 -90
rect 1308 -94 1317 -92
rect 1176 -97 1178 -94
rect 1123 -120 1125 -115
rect 1133 -120 1135 -115
rect 1143 -117 1145 -113
rect 1054 -126 1056 -122
rect 1075 -126 1077 -122
rect 1082 -126 1084 -122
rect 1176 -115 1178 -110
rect 1163 -126 1165 -122
rect 1186 -124 1188 -119
rect 1193 -124 1195 -119
rect 1308 -97 1310 -94
rect 1321 -97 1323 -84
rect 1342 -92 1344 -82
rect 1352 -85 1354 -82
rect 1362 -85 1364 -82
rect 1348 -87 1354 -85
rect 1348 -89 1350 -87
rect 1352 -89 1354 -87
rect 1348 -91 1354 -89
rect 1358 -87 1364 -85
rect 1358 -89 1360 -87
rect 1362 -89 1364 -87
rect 1358 -91 1364 -89
rect 1338 -94 1344 -92
rect 1338 -96 1340 -94
rect 1342 -96 1344 -94
rect 1308 -115 1310 -110
rect 1211 -126 1213 -122
rect 1221 -126 1223 -122
rect 1231 -126 1233 -122
rect 1253 -126 1255 -122
rect 1263 -126 1265 -122
rect 1273 -126 1275 -122
rect 1291 -124 1293 -119
rect 1298 -124 1300 -119
rect 1338 -98 1344 -96
rect 1342 -101 1344 -98
rect 1349 -101 1351 -91
rect 1362 -94 1364 -91
rect 1390 -93 1392 -80
rect 1397 -85 1399 -80
rect 1410 -85 1412 -80
rect 1396 -87 1402 -85
rect 1396 -89 1398 -87
rect 1400 -89 1402 -87
rect 1396 -91 1402 -89
rect 1406 -87 1412 -85
rect 1406 -89 1408 -87
rect 1410 -89 1412 -87
rect 1406 -91 1412 -89
rect 1386 -95 1392 -93
rect 1386 -97 1388 -95
rect 1390 -97 1392 -95
rect 1386 -99 1392 -97
rect 1390 -102 1392 -99
rect 1400 -102 1402 -91
rect 1410 -95 1412 -91
rect 1430 -82 1432 -80
rect 1434 -82 1436 -80
rect 1430 -84 1436 -82
rect 1362 -117 1364 -112
rect 1430 -97 1432 -84
rect 1440 -88 1442 -75
rect 1436 -90 1442 -88
rect 1436 -92 1438 -90
rect 1440 -92 1442 -90
rect 1450 -85 1452 -82
rect 1460 -85 1462 -82
rect 1480 -85 1482 -82
rect 1487 -85 1489 -82
rect 1498 -85 1500 -76
rect 1520 -85 1522 -76
rect 1558 -68 1560 -63
rect 1568 -68 1570 -63
rect 1578 -65 1580 -60
rect 1588 -62 1590 -58
rect 1531 -85 1533 -82
rect 1538 -85 1540 -82
rect 1558 -85 1560 -82
rect 1568 -85 1570 -82
rect 1450 -87 1456 -85
rect 1450 -89 1452 -87
rect 1454 -89 1456 -87
rect 1450 -91 1456 -89
rect 1460 -87 1482 -85
rect 1460 -89 1471 -87
rect 1473 -89 1478 -87
rect 1480 -89 1482 -87
rect 1460 -91 1482 -89
rect 1486 -87 1492 -85
rect 1486 -89 1488 -87
rect 1490 -89 1492 -87
rect 1486 -91 1492 -89
rect 1496 -87 1502 -85
rect 1496 -89 1498 -87
rect 1500 -89 1502 -87
rect 1496 -91 1502 -89
rect 1518 -87 1524 -85
rect 1518 -89 1520 -87
rect 1522 -89 1524 -87
rect 1518 -91 1524 -89
rect 1528 -87 1534 -85
rect 1528 -89 1530 -87
rect 1532 -89 1534 -87
rect 1528 -91 1534 -89
rect 1538 -87 1560 -85
rect 1538 -89 1540 -87
rect 1542 -89 1547 -87
rect 1549 -89 1560 -87
rect 1538 -91 1560 -89
rect 1564 -87 1570 -85
rect 1564 -89 1566 -87
rect 1568 -89 1570 -87
rect 1564 -91 1570 -89
rect 1578 -88 1580 -75
rect 1588 -78 1590 -75
rect 1584 -80 1590 -78
rect 1584 -82 1586 -80
rect 1588 -82 1590 -80
rect 1609 -76 1611 -71
rect 1619 -76 1621 -71
rect 1629 -73 1631 -68
rect 1657 -69 1659 -64
rect 1664 -69 1666 -64
rect 1697 -62 1699 -58
rect 1677 -71 1679 -67
rect 1707 -65 1709 -60
rect 1747 -62 1749 -58
rect 1754 -62 1756 -58
rect 1765 -62 1767 -58
rect 1787 -62 1789 -58
rect 1798 -62 1800 -58
rect 1805 -62 1807 -58
rect 1717 -68 1719 -63
rect 1727 -68 1729 -63
rect 1697 -78 1699 -75
rect 1697 -80 1703 -78
rect 1584 -84 1590 -82
rect 1578 -90 1584 -88
rect 1436 -94 1445 -92
rect 1453 -94 1455 -91
rect 1460 -94 1462 -91
rect 1478 -94 1480 -91
rect 1488 -94 1490 -91
rect 1498 -94 1500 -91
rect 1520 -94 1522 -91
rect 1530 -94 1532 -91
rect 1540 -94 1542 -91
rect 1558 -94 1560 -91
rect 1565 -94 1567 -91
rect 1578 -92 1580 -90
rect 1582 -92 1584 -90
rect 1575 -94 1584 -92
rect 1443 -97 1445 -94
rect 1390 -120 1392 -115
rect 1400 -120 1402 -115
rect 1410 -117 1412 -113
rect 1321 -126 1323 -122
rect 1342 -126 1344 -122
rect 1349 -126 1351 -122
rect 1443 -115 1445 -110
rect 1430 -126 1432 -122
rect 1453 -124 1455 -119
rect 1460 -124 1462 -119
rect 1575 -97 1577 -94
rect 1588 -97 1590 -84
rect 1609 -92 1611 -82
rect 1619 -85 1621 -82
rect 1629 -85 1631 -82
rect 1615 -87 1621 -85
rect 1615 -89 1617 -87
rect 1619 -89 1621 -87
rect 1615 -91 1621 -89
rect 1625 -87 1631 -85
rect 1625 -89 1627 -87
rect 1629 -89 1631 -87
rect 1625 -91 1631 -89
rect 1605 -94 1611 -92
rect 1605 -96 1607 -94
rect 1609 -96 1611 -94
rect 1575 -115 1577 -110
rect 1478 -126 1480 -122
rect 1488 -126 1490 -122
rect 1498 -126 1500 -122
rect 1520 -126 1522 -122
rect 1530 -126 1532 -122
rect 1540 -126 1542 -122
rect 1558 -124 1560 -119
rect 1565 -124 1567 -119
rect 1605 -98 1611 -96
rect 1609 -101 1611 -98
rect 1616 -101 1618 -91
rect 1629 -94 1631 -91
rect 1657 -93 1659 -80
rect 1664 -85 1666 -80
rect 1677 -85 1679 -80
rect 1663 -87 1669 -85
rect 1663 -89 1665 -87
rect 1667 -89 1669 -87
rect 1663 -91 1669 -89
rect 1673 -87 1679 -85
rect 1673 -89 1675 -87
rect 1677 -89 1679 -87
rect 1673 -91 1679 -89
rect 1653 -95 1659 -93
rect 1653 -97 1655 -95
rect 1657 -97 1659 -95
rect 1653 -99 1659 -97
rect 1657 -102 1659 -99
rect 1667 -102 1669 -91
rect 1677 -95 1679 -91
rect 1697 -82 1699 -80
rect 1701 -82 1703 -80
rect 1697 -84 1703 -82
rect 1629 -117 1631 -112
rect 1697 -97 1699 -84
rect 1707 -88 1709 -75
rect 1703 -90 1709 -88
rect 1703 -92 1705 -90
rect 1707 -92 1709 -90
rect 1717 -85 1719 -82
rect 1727 -85 1729 -82
rect 1747 -85 1749 -82
rect 1754 -85 1756 -82
rect 1765 -85 1767 -76
rect 1787 -85 1789 -76
rect 1825 -68 1827 -63
rect 1835 -68 1837 -63
rect 1845 -65 1847 -60
rect 1855 -62 1857 -58
rect 1922 -60 1947 -58
rect 1922 -68 1924 -60
rect 1935 -68 1937 -64
rect 1945 -68 1947 -60
rect 1955 -65 1957 -60
rect 1962 -65 1964 -60
rect 1983 -62 1985 -58
rect 1798 -85 1800 -82
rect 1805 -85 1807 -82
rect 1825 -85 1827 -82
rect 1835 -85 1837 -82
rect 1717 -87 1723 -85
rect 1717 -89 1719 -87
rect 1721 -89 1723 -87
rect 1717 -91 1723 -89
rect 1727 -87 1749 -85
rect 1727 -89 1738 -87
rect 1740 -89 1745 -87
rect 1747 -89 1749 -87
rect 1727 -91 1749 -89
rect 1753 -87 1759 -85
rect 1753 -89 1755 -87
rect 1757 -89 1759 -87
rect 1753 -91 1759 -89
rect 1763 -87 1769 -85
rect 1763 -89 1765 -87
rect 1767 -89 1769 -87
rect 1763 -91 1769 -89
rect 1785 -87 1791 -85
rect 1785 -89 1787 -87
rect 1789 -89 1791 -87
rect 1785 -91 1791 -89
rect 1795 -87 1801 -85
rect 1795 -89 1797 -87
rect 1799 -89 1801 -87
rect 1795 -91 1801 -89
rect 1805 -87 1827 -85
rect 1805 -89 1807 -87
rect 1809 -89 1814 -87
rect 1816 -89 1827 -87
rect 1805 -91 1827 -89
rect 1831 -87 1837 -85
rect 1831 -89 1833 -87
rect 1835 -89 1837 -87
rect 1831 -91 1837 -89
rect 1845 -88 1847 -75
rect 1855 -78 1857 -75
rect 1851 -80 1857 -78
rect 1851 -82 1853 -80
rect 1855 -82 1857 -80
rect 1876 -76 1878 -71
rect 1886 -76 1888 -71
rect 1896 -73 1898 -68
rect 1919 -70 1924 -68
rect 1919 -73 1921 -70
rect 1993 -65 1995 -60
rect 2033 -62 2035 -58
rect 2040 -62 2042 -58
rect 2051 -62 2053 -58
rect 2073 -62 2075 -58
rect 2084 -62 2086 -58
rect 2091 -62 2093 -58
rect 2003 -68 2005 -63
rect 2013 -68 2015 -63
rect 1935 -80 1937 -77
rect 1928 -82 1937 -80
rect 1945 -81 1947 -77
rect 1955 -80 1957 -77
rect 1851 -84 1857 -82
rect 1845 -90 1851 -88
rect 1703 -94 1712 -92
rect 1720 -94 1722 -91
rect 1727 -94 1729 -91
rect 1745 -94 1747 -91
rect 1755 -94 1757 -91
rect 1765 -94 1767 -91
rect 1787 -94 1789 -91
rect 1797 -94 1799 -91
rect 1807 -94 1809 -91
rect 1825 -94 1827 -91
rect 1832 -94 1834 -91
rect 1845 -92 1847 -90
rect 1849 -92 1851 -90
rect 1842 -94 1851 -92
rect 1710 -97 1712 -94
rect 1657 -120 1659 -115
rect 1667 -120 1669 -115
rect 1677 -117 1679 -113
rect 1588 -126 1590 -122
rect 1609 -126 1611 -122
rect 1616 -126 1618 -122
rect 1710 -115 1712 -110
rect 1697 -126 1699 -122
rect 1720 -124 1722 -119
rect 1727 -124 1729 -119
rect 1842 -97 1844 -94
rect 1855 -97 1857 -84
rect 1876 -92 1878 -82
rect 1886 -85 1888 -82
rect 1896 -85 1898 -82
rect 1882 -87 1888 -85
rect 1882 -89 1884 -87
rect 1886 -89 1888 -87
rect 1882 -91 1888 -89
rect 1892 -87 1898 -85
rect 1892 -89 1894 -87
rect 1896 -89 1898 -87
rect 1892 -91 1898 -89
rect 1919 -90 1921 -82
rect 1928 -84 1930 -82
rect 1932 -84 1937 -82
rect 1928 -86 1937 -84
rect 1953 -82 1957 -80
rect 1953 -85 1955 -82
rect 1935 -90 1937 -86
rect 1949 -87 1955 -85
rect 1962 -86 1964 -77
rect 1983 -78 1985 -75
rect 1983 -80 1989 -78
rect 1983 -82 1985 -80
rect 1987 -82 1989 -80
rect 1983 -84 1989 -82
rect 1949 -89 1951 -87
rect 1953 -89 1955 -87
rect 1872 -94 1878 -92
rect 1872 -96 1874 -94
rect 1876 -96 1878 -94
rect 1842 -115 1844 -110
rect 1745 -126 1747 -122
rect 1755 -126 1757 -122
rect 1765 -126 1767 -122
rect 1787 -126 1789 -122
rect 1797 -126 1799 -122
rect 1807 -126 1809 -122
rect 1825 -124 1827 -119
rect 1832 -124 1834 -119
rect 1872 -98 1878 -96
rect 1876 -101 1878 -98
rect 1883 -101 1885 -91
rect 1896 -94 1898 -91
rect 1916 -92 1929 -90
rect 1935 -92 1945 -90
rect 1949 -91 1955 -89
rect 1916 -93 1918 -92
rect 1912 -95 1918 -93
rect 1927 -95 1929 -92
rect 1943 -95 1945 -92
rect 1953 -95 1955 -91
rect 1959 -88 1965 -86
rect 1959 -90 1961 -88
rect 1963 -90 1965 -88
rect 1959 -92 1965 -90
rect 1963 -95 1965 -92
rect 1912 -97 1914 -95
rect 1916 -97 1918 -95
rect 1912 -99 1918 -97
rect 1896 -117 1898 -112
rect 1855 -126 1857 -122
rect 1876 -126 1878 -122
rect 1883 -126 1885 -122
rect 1943 -117 1945 -113
rect 1953 -117 1955 -113
rect 1927 -126 1929 -122
rect 1983 -97 1985 -84
rect 1993 -88 1995 -75
rect 1989 -90 1995 -88
rect 1989 -92 1991 -90
rect 1993 -92 1995 -90
rect 2003 -85 2005 -82
rect 2013 -85 2015 -82
rect 2033 -85 2035 -82
rect 2040 -85 2042 -82
rect 2051 -85 2053 -76
rect 2073 -85 2075 -76
rect 2111 -68 2113 -63
rect 2121 -68 2123 -63
rect 2131 -65 2133 -60
rect 2141 -62 2143 -58
rect 2206 -60 2225 -58
rect 2084 -85 2086 -82
rect 2091 -85 2093 -82
rect 2111 -85 2113 -82
rect 2121 -85 2123 -82
rect 2003 -87 2009 -85
rect 2003 -89 2005 -87
rect 2007 -89 2009 -87
rect 2003 -91 2009 -89
rect 2013 -87 2035 -85
rect 2013 -89 2024 -87
rect 2026 -89 2031 -87
rect 2033 -89 2035 -87
rect 2013 -91 2035 -89
rect 2039 -87 2045 -85
rect 2039 -89 2041 -87
rect 2043 -89 2045 -87
rect 2039 -91 2045 -89
rect 2049 -87 2055 -85
rect 2049 -89 2051 -87
rect 2053 -89 2055 -87
rect 2049 -91 2055 -89
rect 2071 -87 2077 -85
rect 2071 -89 2073 -87
rect 2075 -89 2077 -87
rect 2071 -91 2077 -89
rect 2081 -87 2087 -85
rect 2081 -89 2083 -87
rect 2085 -89 2087 -87
rect 2081 -91 2087 -89
rect 2091 -87 2113 -85
rect 2091 -89 2093 -87
rect 2095 -89 2100 -87
rect 2102 -89 2113 -87
rect 2091 -91 2113 -89
rect 2117 -87 2123 -85
rect 2117 -89 2119 -87
rect 2121 -89 2123 -87
rect 2117 -91 2123 -89
rect 2131 -88 2133 -75
rect 2141 -78 2143 -75
rect 2137 -80 2143 -78
rect 2137 -82 2139 -80
rect 2141 -82 2143 -80
rect 2162 -76 2164 -71
rect 2172 -76 2174 -71
rect 2182 -73 2184 -68
rect 2206 -70 2208 -60
rect 2216 -68 2218 -64
rect 2223 -68 2225 -60
rect 2274 -60 2293 -58
rect 2233 -68 2235 -63
rect 2240 -68 2242 -63
rect 2250 -68 2252 -63
rect 2137 -84 2143 -82
rect 2131 -90 2137 -88
rect 1989 -94 1998 -92
rect 2006 -94 2008 -91
rect 2013 -94 2015 -91
rect 2031 -94 2033 -91
rect 2041 -94 2043 -91
rect 2051 -94 2053 -91
rect 2073 -94 2075 -91
rect 2083 -94 2085 -91
rect 2093 -94 2095 -91
rect 2111 -94 2113 -91
rect 2118 -94 2120 -91
rect 2131 -92 2133 -90
rect 2135 -92 2137 -90
rect 2128 -94 2137 -92
rect 1996 -97 1998 -94
rect 1996 -115 1998 -110
rect 1963 -126 1965 -122
rect 1983 -126 1985 -122
rect 2006 -124 2008 -119
rect 2013 -124 2015 -119
rect 2128 -97 2130 -94
rect 2141 -97 2143 -84
rect 2162 -92 2164 -82
rect 2172 -85 2174 -82
rect 2182 -85 2184 -82
rect 2168 -87 2174 -85
rect 2168 -89 2170 -87
rect 2172 -89 2174 -87
rect 2168 -91 2174 -89
rect 2178 -87 2184 -85
rect 2178 -89 2180 -87
rect 2182 -89 2184 -87
rect 2178 -91 2184 -89
rect 2158 -94 2164 -92
rect 2158 -96 2160 -94
rect 2162 -96 2164 -94
rect 2128 -115 2130 -110
rect 2031 -126 2033 -122
rect 2041 -126 2043 -122
rect 2051 -126 2053 -122
rect 2073 -126 2075 -122
rect 2083 -126 2085 -122
rect 2093 -126 2095 -122
rect 2111 -124 2113 -119
rect 2118 -124 2120 -119
rect 2158 -98 2164 -96
rect 2162 -101 2164 -98
rect 2169 -101 2171 -91
rect 2182 -94 2184 -91
rect 2206 -94 2208 -76
rect 2216 -85 2218 -76
rect 2212 -87 2218 -85
rect 2212 -89 2214 -87
rect 2216 -89 2218 -87
rect 2212 -91 2218 -89
rect 2223 -89 2225 -76
rect 2233 -79 2235 -76
rect 2229 -81 2235 -79
rect 2229 -83 2231 -81
rect 2233 -83 2235 -81
rect 2229 -85 2235 -83
rect 2223 -91 2235 -89
rect 2240 -90 2242 -76
rect 2274 -70 2276 -60
rect 2284 -68 2286 -64
rect 2291 -68 2293 -60
rect 2301 -68 2303 -63
rect 2308 -68 2310 -63
rect 2318 -68 2320 -63
rect 2250 -80 2252 -77
rect 2247 -82 2253 -80
rect 2247 -84 2249 -82
rect 2251 -84 2253 -82
rect 2247 -86 2253 -84
rect 2206 -105 2208 -102
rect 2199 -107 2208 -105
rect 2216 -106 2218 -91
rect 2222 -97 2228 -95
rect 2222 -99 2224 -97
rect 2226 -99 2228 -97
rect 2222 -101 2228 -99
rect 2223 -106 2225 -101
rect 2233 -106 2235 -91
rect 2239 -92 2245 -90
rect 2239 -94 2241 -92
rect 2243 -94 2245 -92
rect 2239 -96 2245 -94
rect 2240 -106 2242 -96
rect 2250 -104 2252 -86
rect 2274 -94 2276 -76
rect 2284 -85 2286 -76
rect 2280 -87 2286 -85
rect 2280 -89 2282 -87
rect 2284 -89 2286 -87
rect 2280 -91 2286 -89
rect 2291 -89 2293 -76
rect 2301 -79 2303 -76
rect 2297 -81 2303 -79
rect 2297 -83 2299 -81
rect 2301 -83 2303 -81
rect 2297 -85 2303 -83
rect 2291 -91 2303 -89
rect 2308 -90 2310 -76
rect 2318 -80 2320 -77
rect 2315 -82 2321 -80
rect 2315 -84 2317 -82
rect 2319 -84 2321 -82
rect 2315 -86 2321 -84
rect 2199 -109 2201 -107
rect 2203 -109 2205 -107
rect 2199 -111 2205 -109
rect 2182 -117 2184 -112
rect 2141 -126 2143 -122
rect 2162 -126 2164 -122
rect 2169 -126 2171 -122
rect 2274 -105 2276 -102
rect 2267 -107 2276 -105
rect 2284 -106 2286 -91
rect 2290 -97 2296 -95
rect 2290 -99 2292 -97
rect 2294 -99 2296 -97
rect 2290 -101 2296 -99
rect 2291 -106 2293 -101
rect 2301 -106 2303 -91
rect 2307 -92 2313 -90
rect 2307 -94 2309 -92
rect 2311 -94 2313 -92
rect 2307 -96 2313 -94
rect 2308 -106 2310 -96
rect 2318 -104 2320 -86
rect 2267 -109 2269 -107
rect 2271 -109 2273 -107
rect 2267 -111 2273 -109
rect 2216 -126 2218 -122
rect 2223 -126 2225 -122
rect 2233 -126 2235 -122
rect 2240 -126 2242 -122
rect 2250 -126 2252 -122
rect 2284 -126 2286 -122
rect 2291 -126 2293 -122
rect 2301 -126 2303 -122
rect 2308 -126 2310 -122
rect 2318 -126 2320 -122
rect 15 -141 17 -136
rect 25 -141 27 -136
rect 95 -134 97 -130
rect 35 -143 37 -139
rect 55 -141 57 -136
rect 65 -141 67 -136
rect 15 -157 17 -154
rect 11 -159 17 -157
rect 11 -161 13 -159
rect 15 -161 17 -159
rect 11 -163 17 -161
rect 15 -176 17 -163
rect 25 -165 27 -154
rect 75 -143 77 -139
rect 55 -157 57 -154
rect 51 -159 57 -157
rect 51 -161 53 -159
rect 55 -161 57 -159
rect 35 -165 37 -161
rect 51 -163 57 -161
rect 21 -167 27 -165
rect 21 -169 23 -167
rect 25 -169 27 -167
rect 21 -171 27 -169
rect 31 -167 37 -165
rect 31 -169 33 -167
rect 35 -169 37 -167
rect 31 -171 37 -169
rect 22 -176 24 -171
rect 35 -176 37 -171
rect 55 -176 57 -163
rect 65 -165 67 -154
rect 118 -137 120 -132
rect 125 -137 127 -132
rect 143 -134 145 -130
rect 153 -134 155 -130
rect 163 -134 165 -130
rect 185 -134 187 -130
rect 195 -134 197 -130
rect 205 -134 207 -130
rect 108 -146 110 -141
rect 75 -165 77 -161
rect 61 -167 67 -165
rect 61 -169 63 -167
rect 65 -169 67 -167
rect 61 -171 67 -169
rect 71 -167 77 -165
rect 71 -169 73 -167
rect 75 -169 77 -167
rect 71 -171 77 -169
rect 62 -176 64 -171
rect 75 -176 77 -171
rect 95 -172 97 -159
rect 108 -162 110 -159
rect 223 -137 225 -132
rect 230 -137 232 -132
rect 253 -134 255 -130
rect 274 -134 276 -130
rect 281 -134 283 -130
rect 240 -146 242 -141
rect 362 -134 364 -130
rect 294 -144 296 -139
rect 322 -141 324 -136
rect 332 -141 334 -136
rect 274 -158 276 -155
rect 240 -162 242 -159
rect 101 -164 110 -162
rect 101 -166 103 -164
rect 105 -166 107 -164
rect 118 -165 120 -162
rect 125 -165 127 -162
rect 143 -165 145 -162
rect 153 -165 155 -162
rect 163 -165 165 -162
rect 185 -165 187 -162
rect 195 -165 197 -162
rect 205 -165 207 -162
rect 223 -165 225 -162
rect 230 -165 232 -162
rect 240 -164 249 -162
rect 101 -168 107 -166
rect 95 -174 101 -172
rect 95 -176 97 -174
rect 99 -176 101 -174
rect 15 -192 17 -187
rect 22 -192 24 -187
rect 35 -189 37 -185
rect 95 -178 101 -176
rect 95 -181 97 -178
rect 105 -181 107 -168
rect 115 -167 121 -165
rect 115 -169 117 -167
rect 119 -169 121 -167
rect 115 -171 121 -169
rect 125 -167 147 -165
rect 125 -169 136 -167
rect 138 -169 143 -167
rect 145 -169 147 -167
rect 125 -171 147 -169
rect 151 -167 157 -165
rect 151 -169 153 -167
rect 155 -169 157 -167
rect 151 -171 157 -169
rect 161 -167 167 -165
rect 161 -169 163 -167
rect 165 -169 167 -167
rect 161 -171 167 -169
rect 183 -167 189 -165
rect 183 -169 185 -167
rect 187 -169 189 -167
rect 183 -171 189 -169
rect 193 -167 199 -165
rect 193 -169 195 -167
rect 197 -169 199 -167
rect 193 -171 199 -169
rect 203 -167 225 -165
rect 203 -169 205 -167
rect 207 -169 212 -167
rect 214 -169 225 -167
rect 203 -171 225 -169
rect 229 -167 235 -165
rect 229 -169 231 -167
rect 233 -169 235 -167
rect 229 -171 235 -169
rect 115 -174 117 -171
rect 125 -174 127 -171
rect 145 -174 147 -171
rect 152 -174 154 -171
rect 55 -192 57 -187
rect 62 -192 64 -187
rect 75 -189 77 -185
rect 95 -198 97 -194
rect 105 -196 107 -191
rect 115 -193 117 -188
rect 125 -193 127 -188
rect 163 -180 165 -171
rect 185 -180 187 -171
rect 196 -174 198 -171
rect 203 -174 205 -171
rect 223 -174 225 -171
rect 233 -174 235 -171
rect 243 -166 245 -164
rect 247 -166 249 -164
rect 243 -168 249 -166
rect 243 -181 245 -168
rect 253 -172 255 -159
rect 270 -160 276 -158
rect 270 -162 272 -160
rect 274 -162 276 -160
rect 270 -164 276 -162
rect 249 -174 255 -172
rect 274 -174 276 -164
rect 281 -165 283 -155
rect 342 -143 344 -139
rect 322 -157 324 -154
rect 318 -159 324 -157
rect 318 -161 320 -159
rect 322 -161 324 -159
rect 294 -165 296 -162
rect 318 -163 324 -161
rect 280 -167 286 -165
rect 280 -169 282 -167
rect 284 -169 286 -167
rect 280 -171 286 -169
rect 290 -167 296 -165
rect 290 -169 292 -167
rect 294 -169 296 -167
rect 290 -171 296 -169
rect 284 -174 286 -171
rect 294 -174 296 -171
rect 249 -176 251 -174
rect 253 -176 255 -174
rect 249 -178 255 -176
rect 253 -181 255 -178
rect 223 -193 225 -188
rect 233 -193 235 -188
rect 145 -198 147 -194
rect 152 -198 154 -194
rect 163 -198 165 -194
rect 185 -198 187 -194
rect 196 -198 198 -194
rect 203 -198 205 -194
rect 243 -196 245 -191
rect 274 -185 276 -180
rect 284 -185 286 -180
rect 322 -176 324 -163
rect 332 -165 334 -154
rect 385 -137 387 -132
rect 392 -137 394 -132
rect 410 -134 412 -130
rect 420 -134 422 -130
rect 430 -134 432 -130
rect 452 -134 454 -130
rect 462 -134 464 -130
rect 472 -134 474 -130
rect 375 -146 377 -141
rect 342 -165 344 -161
rect 328 -167 334 -165
rect 328 -169 330 -167
rect 332 -169 334 -167
rect 328 -171 334 -169
rect 338 -167 344 -165
rect 338 -169 340 -167
rect 342 -169 344 -167
rect 338 -171 344 -169
rect 329 -176 331 -171
rect 342 -176 344 -171
rect 362 -172 364 -159
rect 375 -162 377 -159
rect 490 -137 492 -132
rect 497 -137 499 -132
rect 520 -134 522 -130
rect 541 -134 543 -130
rect 548 -134 550 -130
rect 507 -146 509 -141
rect 629 -134 631 -130
rect 561 -144 563 -139
rect 589 -141 591 -136
rect 599 -141 601 -136
rect 541 -158 543 -155
rect 507 -162 509 -159
rect 368 -164 377 -162
rect 368 -166 370 -164
rect 372 -166 374 -164
rect 385 -165 387 -162
rect 392 -165 394 -162
rect 410 -165 412 -162
rect 420 -165 422 -162
rect 430 -165 432 -162
rect 452 -165 454 -162
rect 462 -165 464 -162
rect 472 -165 474 -162
rect 490 -165 492 -162
rect 497 -165 499 -162
rect 507 -164 516 -162
rect 368 -168 374 -166
rect 362 -174 368 -172
rect 362 -176 364 -174
rect 366 -176 368 -174
rect 294 -188 296 -183
rect 362 -178 368 -176
rect 362 -181 364 -178
rect 372 -181 374 -168
rect 382 -167 388 -165
rect 382 -169 384 -167
rect 386 -169 388 -167
rect 382 -171 388 -169
rect 392 -167 414 -165
rect 392 -169 403 -167
rect 405 -169 410 -167
rect 412 -169 414 -167
rect 392 -171 414 -169
rect 418 -167 424 -165
rect 418 -169 420 -167
rect 422 -169 424 -167
rect 418 -171 424 -169
rect 428 -167 434 -165
rect 428 -169 430 -167
rect 432 -169 434 -167
rect 428 -171 434 -169
rect 450 -167 456 -165
rect 450 -169 452 -167
rect 454 -169 456 -167
rect 450 -171 456 -169
rect 460 -167 466 -165
rect 460 -169 462 -167
rect 464 -169 466 -167
rect 460 -171 466 -169
rect 470 -167 492 -165
rect 470 -169 472 -167
rect 474 -169 479 -167
rect 481 -169 492 -167
rect 470 -171 492 -169
rect 496 -167 502 -165
rect 496 -169 498 -167
rect 500 -169 502 -167
rect 496 -171 502 -169
rect 382 -174 384 -171
rect 392 -174 394 -171
rect 412 -174 414 -171
rect 419 -174 421 -171
rect 322 -192 324 -187
rect 329 -192 331 -187
rect 253 -198 255 -194
rect 342 -189 344 -185
rect 362 -198 364 -194
rect 372 -196 374 -191
rect 382 -193 384 -188
rect 392 -193 394 -188
rect 430 -180 432 -171
rect 452 -180 454 -171
rect 463 -174 465 -171
rect 470 -174 472 -171
rect 490 -174 492 -171
rect 500 -174 502 -171
rect 510 -166 512 -164
rect 514 -166 516 -164
rect 510 -168 516 -166
rect 510 -181 512 -168
rect 520 -172 522 -159
rect 537 -160 543 -158
rect 537 -162 539 -160
rect 541 -162 543 -160
rect 537 -164 543 -162
rect 516 -174 522 -172
rect 541 -174 543 -164
rect 548 -165 550 -155
rect 609 -143 611 -139
rect 589 -157 591 -154
rect 585 -159 591 -157
rect 585 -161 587 -159
rect 589 -161 591 -159
rect 561 -165 563 -162
rect 585 -163 591 -161
rect 547 -167 553 -165
rect 547 -169 549 -167
rect 551 -169 553 -167
rect 547 -171 553 -169
rect 557 -167 563 -165
rect 557 -169 559 -167
rect 561 -169 563 -167
rect 557 -171 563 -169
rect 551 -174 553 -171
rect 561 -174 563 -171
rect 516 -176 518 -174
rect 520 -176 522 -174
rect 516 -178 522 -176
rect 520 -181 522 -178
rect 490 -193 492 -188
rect 500 -193 502 -188
rect 412 -198 414 -194
rect 419 -198 421 -194
rect 430 -198 432 -194
rect 452 -198 454 -194
rect 463 -198 465 -194
rect 470 -198 472 -194
rect 510 -196 512 -191
rect 541 -185 543 -180
rect 551 -185 553 -180
rect 589 -176 591 -163
rect 599 -165 601 -154
rect 652 -137 654 -132
rect 659 -137 661 -132
rect 677 -134 679 -130
rect 687 -134 689 -130
rect 697 -134 699 -130
rect 719 -134 721 -130
rect 729 -134 731 -130
rect 739 -134 741 -130
rect 642 -146 644 -141
rect 609 -165 611 -161
rect 595 -167 601 -165
rect 595 -169 597 -167
rect 599 -169 601 -167
rect 595 -171 601 -169
rect 605 -167 611 -165
rect 605 -169 607 -167
rect 609 -169 611 -167
rect 605 -171 611 -169
rect 596 -176 598 -171
rect 609 -176 611 -171
rect 629 -172 631 -159
rect 642 -162 644 -159
rect 757 -137 759 -132
rect 764 -137 766 -132
rect 787 -134 789 -130
rect 808 -134 810 -130
rect 815 -134 817 -130
rect 774 -146 776 -141
rect 896 -134 898 -130
rect 828 -144 830 -139
rect 856 -141 858 -136
rect 866 -141 868 -136
rect 808 -158 810 -155
rect 774 -162 776 -159
rect 635 -164 644 -162
rect 635 -166 637 -164
rect 639 -166 641 -164
rect 652 -165 654 -162
rect 659 -165 661 -162
rect 677 -165 679 -162
rect 687 -165 689 -162
rect 697 -165 699 -162
rect 719 -165 721 -162
rect 729 -165 731 -162
rect 739 -165 741 -162
rect 757 -165 759 -162
rect 764 -165 766 -162
rect 774 -164 783 -162
rect 635 -168 641 -166
rect 629 -174 635 -172
rect 629 -176 631 -174
rect 633 -176 635 -174
rect 561 -188 563 -183
rect 629 -178 635 -176
rect 629 -181 631 -178
rect 639 -181 641 -168
rect 649 -167 655 -165
rect 649 -169 651 -167
rect 653 -169 655 -167
rect 649 -171 655 -169
rect 659 -167 681 -165
rect 659 -169 670 -167
rect 672 -169 677 -167
rect 679 -169 681 -167
rect 659 -171 681 -169
rect 685 -167 691 -165
rect 685 -169 687 -167
rect 689 -169 691 -167
rect 685 -171 691 -169
rect 695 -167 701 -165
rect 695 -169 697 -167
rect 699 -169 701 -167
rect 695 -171 701 -169
rect 717 -167 723 -165
rect 717 -169 719 -167
rect 721 -169 723 -167
rect 717 -171 723 -169
rect 727 -167 733 -165
rect 727 -169 729 -167
rect 731 -169 733 -167
rect 727 -171 733 -169
rect 737 -167 759 -165
rect 737 -169 739 -167
rect 741 -169 746 -167
rect 748 -169 759 -167
rect 737 -171 759 -169
rect 763 -167 769 -165
rect 763 -169 765 -167
rect 767 -169 769 -167
rect 763 -171 769 -169
rect 649 -174 651 -171
rect 659 -174 661 -171
rect 679 -174 681 -171
rect 686 -174 688 -171
rect 589 -192 591 -187
rect 596 -192 598 -187
rect 520 -198 522 -194
rect 609 -189 611 -185
rect 629 -198 631 -194
rect 639 -196 641 -191
rect 649 -193 651 -188
rect 659 -193 661 -188
rect 697 -180 699 -171
rect 719 -180 721 -171
rect 730 -174 732 -171
rect 737 -174 739 -171
rect 757 -174 759 -171
rect 767 -174 769 -171
rect 777 -166 779 -164
rect 781 -166 783 -164
rect 777 -168 783 -166
rect 777 -181 779 -168
rect 787 -172 789 -159
rect 804 -160 810 -158
rect 804 -162 806 -160
rect 808 -162 810 -160
rect 804 -164 810 -162
rect 783 -174 789 -172
rect 808 -174 810 -164
rect 815 -165 817 -155
rect 876 -143 878 -139
rect 856 -157 858 -154
rect 852 -159 858 -157
rect 852 -161 854 -159
rect 856 -161 858 -159
rect 828 -165 830 -162
rect 852 -163 858 -161
rect 814 -167 820 -165
rect 814 -169 816 -167
rect 818 -169 820 -167
rect 814 -171 820 -169
rect 824 -167 830 -165
rect 824 -169 826 -167
rect 828 -169 830 -167
rect 824 -171 830 -169
rect 818 -174 820 -171
rect 828 -174 830 -171
rect 783 -176 785 -174
rect 787 -176 789 -174
rect 783 -178 789 -176
rect 787 -181 789 -178
rect 757 -193 759 -188
rect 767 -193 769 -188
rect 679 -198 681 -194
rect 686 -198 688 -194
rect 697 -198 699 -194
rect 719 -198 721 -194
rect 730 -198 732 -194
rect 737 -198 739 -194
rect 777 -196 779 -191
rect 808 -185 810 -180
rect 818 -185 820 -180
rect 856 -176 858 -163
rect 866 -165 868 -154
rect 919 -137 921 -132
rect 926 -137 928 -132
rect 944 -134 946 -130
rect 954 -134 956 -130
rect 964 -134 966 -130
rect 986 -134 988 -130
rect 996 -134 998 -130
rect 1006 -134 1008 -130
rect 909 -146 911 -141
rect 876 -165 878 -161
rect 862 -167 868 -165
rect 862 -169 864 -167
rect 866 -169 868 -167
rect 862 -171 868 -169
rect 872 -167 878 -165
rect 872 -169 874 -167
rect 876 -169 878 -167
rect 872 -171 878 -169
rect 863 -176 865 -171
rect 876 -176 878 -171
rect 896 -172 898 -159
rect 909 -162 911 -159
rect 1024 -137 1026 -132
rect 1031 -137 1033 -132
rect 1054 -134 1056 -130
rect 1075 -134 1077 -130
rect 1082 -134 1084 -130
rect 1041 -146 1043 -141
rect 1163 -134 1165 -130
rect 1095 -144 1097 -139
rect 1123 -141 1125 -136
rect 1133 -141 1135 -136
rect 1075 -158 1077 -155
rect 1041 -162 1043 -159
rect 902 -164 911 -162
rect 902 -166 904 -164
rect 906 -166 908 -164
rect 919 -165 921 -162
rect 926 -165 928 -162
rect 944 -165 946 -162
rect 954 -165 956 -162
rect 964 -165 966 -162
rect 986 -165 988 -162
rect 996 -165 998 -162
rect 1006 -165 1008 -162
rect 1024 -165 1026 -162
rect 1031 -165 1033 -162
rect 1041 -164 1050 -162
rect 902 -168 908 -166
rect 896 -174 902 -172
rect 896 -176 898 -174
rect 900 -176 902 -174
rect 828 -188 830 -183
rect 896 -178 902 -176
rect 896 -181 898 -178
rect 906 -181 908 -168
rect 916 -167 922 -165
rect 916 -169 918 -167
rect 920 -169 922 -167
rect 916 -171 922 -169
rect 926 -167 948 -165
rect 926 -169 937 -167
rect 939 -169 944 -167
rect 946 -169 948 -167
rect 926 -171 948 -169
rect 952 -167 958 -165
rect 952 -169 954 -167
rect 956 -169 958 -167
rect 952 -171 958 -169
rect 962 -167 968 -165
rect 962 -169 964 -167
rect 966 -169 968 -167
rect 962 -171 968 -169
rect 984 -167 990 -165
rect 984 -169 986 -167
rect 988 -169 990 -167
rect 984 -171 990 -169
rect 994 -167 1000 -165
rect 994 -169 996 -167
rect 998 -169 1000 -167
rect 994 -171 1000 -169
rect 1004 -167 1026 -165
rect 1004 -169 1006 -167
rect 1008 -169 1013 -167
rect 1015 -169 1026 -167
rect 1004 -171 1026 -169
rect 1030 -167 1036 -165
rect 1030 -169 1032 -167
rect 1034 -169 1036 -167
rect 1030 -171 1036 -169
rect 916 -174 918 -171
rect 926 -174 928 -171
rect 946 -174 948 -171
rect 953 -174 955 -171
rect 856 -192 858 -187
rect 863 -192 865 -187
rect 787 -198 789 -194
rect 876 -189 878 -185
rect 896 -198 898 -194
rect 906 -196 908 -191
rect 916 -193 918 -188
rect 926 -193 928 -188
rect 964 -180 966 -171
rect 986 -180 988 -171
rect 997 -174 999 -171
rect 1004 -174 1006 -171
rect 1024 -174 1026 -171
rect 1034 -174 1036 -171
rect 1044 -166 1046 -164
rect 1048 -166 1050 -164
rect 1044 -168 1050 -166
rect 1044 -181 1046 -168
rect 1054 -172 1056 -159
rect 1071 -160 1077 -158
rect 1071 -162 1073 -160
rect 1075 -162 1077 -160
rect 1071 -164 1077 -162
rect 1050 -174 1056 -172
rect 1075 -174 1077 -164
rect 1082 -165 1084 -155
rect 1143 -143 1145 -139
rect 1123 -157 1125 -154
rect 1119 -159 1125 -157
rect 1119 -161 1121 -159
rect 1123 -161 1125 -159
rect 1095 -165 1097 -162
rect 1119 -163 1125 -161
rect 1081 -167 1087 -165
rect 1081 -169 1083 -167
rect 1085 -169 1087 -167
rect 1081 -171 1087 -169
rect 1091 -167 1097 -165
rect 1091 -169 1093 -167
rect 1095 -169 1097 -167
rect 1091 -171 1097 -169
rect 1085 -174 1087 -171
rect 1095 -174 1097 -171
rect 1050 -176 1052 -174
rect 1054 -176 1056 -174
rect 1050 -178 1056 -176
rect 1054 -181 1056 -178
rect 1024 -193 1026 -188
rect 1034 -193 1036 -188
rect 946 -198 948 -194
rect 953 -198 955 -194
rect 964 -198 966 -194
rect 986 -198 988 -194
rect 997 -198 999 -194
rect 1004 -198 1006 -194
rect 1044 -196 1046 -191
rect 1075 -185 1077 -180
rect 1085 -185 1087 -180
rect 1123 -176 1125 -163
rect 1133 -165 1135 -154
rect 1186 -137 1188 -132
rect 1193 -137 1195 -132
rect 1211 -134 1213 -130
rect 1221 -134 1223 -130
rect 1231 -134 1233 -130
rect 1253 -134 1255 -130
rect 1263 -134 1265 -130
rect 1273 -134 1275 -130
rect 1176 -146 1178 -141
rect 1143 -165 1145 -161
rect 1129 -167 1135 -165
rect 1129 -169 1131 -167
rect 1133 -169 1135 -167
rect 1129 -171 1135 -169
rect 1139 -167 1145 -165
rect 1139 -169 1141 -167
rect 1143 -169 1145 -167
rect 1139 -171 1145 -169
rect 1130 -176 1132 -171
rect 1143 -176 1145 -171
rect 1163 -172 1165 -159
rect 1176 -162 1178 -159
rect 1291 -137 1293 -132
rect 1298 -137 1300 -132
rect 1321 -134 1323 -130
rect 1342 -134 1344 -130
rect 1349 -134 1351 -130
rect 1308 -146 1310 -141
rect 1430 -134 1432 -130
rect 1362 -144 1364 -139
rect 1390 -141 1392 -136
rect 1400 -141 1402 -136
rect 1342 -158 1344 -155
rect 1308 -162 1310 -159
rect 1169 -164 1178 -162
rect 1169 -166 1171 -164
rect 1173 -166 1175 -164
rect 1186 -165 1188 -162
rect 1193 -165 1195 -162
rect 1211 -165 1213 -162
rect 1221 -165 1223 -162
rect 1231 -165 1233 -162
rect 1253 -165 1255 -162
rect 1263 -165 1265 -162
rect 1273 -165 1275 -162
rect 1291 -165 1293 -162
rect 1298 -165 1300 -162
rect 1308 -164 1317 -162
rect 1169 -168 1175 -166
rect 1163 -174 1169 -172
rect 1163 -176 1165 -174
rect 1167 -176 1169 -174
rect 1095 -188 1097 -183
rect 1163 -178 1169 -176
rect 1163 -181 1165 -178
rect 1173 -181 1175 -168
rect 1183 -167 1189 -165
rect 1183 -169 1185 -167
rect 1187 -169 1189 -167
rect 1183 -171 1189 -169
rect 1193 -167 1215 -165
rect 1193 -169 1204 -167
rect 1206 -169 1211 -167
rect 1213 -169 1215 -167
rect 1193 -171 1215 -169
rect 1219 -167 1225 -165
rect 1219 -169 1221 -167
rect 1223 -169 1225 -167
rect 1219 -171 1225 -169
rect 1229 -167 1235 -165
rect 1229 -169 1231 -167
rect 1233 -169 1235 -167
rect 1229 -171 1235 -169
rect 1251 -167 1257 -165
rect 1251 -169 1253 -167
rect 1255 -169 1257 -167
rect 1251 -171 1257 -169
rect 1261 -167 1267 -165
rect 1261 -169 1263 -167
rect 1265 -169 1267 -167
rect 1261 -171 1267 -169
rect 1271 -167 1293 -165
rect 1271 -169 1273 -167
rect 1275 -169 1280 -167
rect 1282 -169 1293 -167
rect 1271 -171 1293 -169
rect 1297 -167 1303 -165
rect 1297 -169 1299 -167
rect 1301 -169 1303 -167
rect 1297 -171 1303 -169
rect 1183 -174 1185 -171
rect 1193 -174 1195 -171
rect 1213 -174 1215 -171
rect 1220 -174 1222 -171
rect 1123 -192 1125 -187
rect 1130 -192 1132 -187
rect 1054 -198 1056 -194
rect 1143 -189 1145 -185
rect 1163 -198 1165 -194
rect 1173 -196 1175 -191
rect 1183 -193 1185 -188
rect 1193 -193 1195 -188
rect 1231 -180 1233 -171
rect 1253 -180 1255 -171
rect 1264 -174 1266 -171
rect 1271 -174 1273 -171
rect 1291 -174 1293 -171
rect 1301 -174 1303 -171
rect 1311 -166 1313 -164
rect 1315 -166 1317 -164
rect 1311 -168 1317 -166
rect 1311 -181 1313 -168
rect 1321 -172 1323 -159
rect 1338 -160 1344 -158
rect 1338 -162 1340 -160
rect 1342 -162 1344 -160
rect 1338 -164 1344 -162
rect 1317 -174 1323 -172
rect 1342 -174 1344 -164
rect 1349 -165 1351 -155
rect 1410 -143 1412 -139
rect 1390 -157 1392 -154
rect 1386 -159 1392 -157
rect 1386 -161 1388 -159
rect 1390 -161 1392 -159
rect 1362 -165 1364 -162
rect 1386 -163 1392 -161
rect 1348 -167 1354 -165
rect 1348 -169 1350 -167
rect 1352 -169 1354 -167
rect 1348 -171 1354 -169
rect 1358 -167 1364 -165
rect 1358 -169 1360 -167
rect 1362 -169 1364 -167
rect 1358 -171 1364 -169
rect 1352 -174 1354 -171
rect 1362 -174 1364 -171
rect 1317 -176 1319 -174
rect 1321 -176 1323 -174
rect 1317 -178 1323 -176
rect 1321 -181 1323 -178
rect 1291 -193 1293 -188
rect 1301 -193 1303 -188
rect 1213 -198 1215 -194
rect 1220 -198 1222 -194
rect 1231 -198 1233 -194
rect 1253 -198 1255 -194
rect 1264 -198 1266 -194
rect 1271 -198 1273 -194
rect 1311 -196 1313 -191
rect 1342 -185 1344 -180
rect 1352 -185 1354 -180
rect 1390 -176 1392 -163
rect 1400 -165 1402 -154
rect 1453 -137 1455 -132
rect 1460 -137 1462 -132
rect 1478 -134 1480 -130
rect 1488 -134 1490 -130
rect 1498 -134 1500 -130
rect 1520 -134 1522 -130
rect 1530 -134 1532 -130
rect 1540 -134 1542 -130
rect 1443 -146 1445 -141
rect 1410 -165 1412 -161
rect 1396 -167 1402 -165
rect 1396 -169 1398 -167
rect 1400 -169 1402 -167
rect 1396 -171 1402 -169
rect 1406 -167 1412 -165
rect 1406 -169 1408 -167
rect 1410 -169 1412 -167
rect 1406 -171 1412 -169
rect 1397 -176 1399 -171
rect 1410 -176 1412 -171
rect 1430 -172 1432 -159
rect 1443 -162 1445 -159
rect 1558 -137 1560 -132
rect 1565 -137 1567 -132
rect 1588 -134 1590 -130
rect 1609 -134 1611 -130
rect 1616 -134 1618 -130
rect 1575 -146 1577 -141
rect 1697 -134 1699 -130
rect 1629 -144 1631 -139
rect 1657 -141 1659 -136
rect 1667 -141 1669 -136
rect 1609 -158 1611 -155
rect 1575 -162 1577 -159
rect 1436 -164 1445 -162
rect 1436 -166 1438 -164
rect 1440 -166 1442 -164
rect 1453 -165 1455 -162
rect 1460 -165 1462 -162
rect 1478 -165 1480 -162
rect 1488 -165 1490 -162
rect 1498 -165 1500 -162
rect 1520 -165 1522 -162
rect 1530 -165 1532 -162
rect 1540 -165 1542 -162
rect 1558 -165 1560 -162
rect 1565 -165 1567 -162
rect 1575 -164 1584 -162
rect 1436 -168 1442 -166
rect 1430 -174 1436 -172
rect 1430 -176 1432 -174
rect 1434 -176 1436 -174
rect 1362 -188 1364 -183
rect 1430 -178 1436 -176
rect 1430 -181 1432 -178
rect 1440 -181 1442 -168
rect 1450 -167 1456 -165
rect 1450 -169 1452 -167
rect 1454 -169 1456 -167
rect 1450 -171 1456 -169
rect 1460 -167 1482 -165
rect 1460 -169 1471 -167
rect 1473 -169 1478 -167
rect 1480 -169 1482 -167
rect 1460 -171 1482 -169
rect 1486 -167 1492 -165
rect 1486 -169 1488 -167
rect 1490 -169 1492 -167
rect 1486 -171 1492 -169
rect 1496 -167 1502 -165
rect 1496 -169 1498 -167
rect 1500 -169 1502 -167
rect 1496 -171 1502 -169
rect 1518 -167 1524 -165
rect 1518 -169 1520 -167
rect 1522 -169 1524 -167
rect 1518 -171 1524 -169
rect 1528 -167 1534 -165
rect 1528 -169 1530 -167
rect 1532 -169 1534 -167
rect 1528 -171 1534 -169
rect 1538 -167 1560 -165
rect 1538 -169 1540 -167
rect 1542 -169 1547 -167
rect 1549 -169 1560 -167
rect 1538 -171 1560 -169
rect 1564 -167 1570 -165
rect 1564 -169 1566 -167
rect 1568 -169 1570 -167
rect 1564 -171 1570 -169
rect 1450 -174 1452 -171
rect 1460 -174 1462 -171
rect 1480 -174 1482 -171
rect 1487 -174 1489 -171
rect 1390 -192 1392 -187
rect 1397 -192 1399 -187
rect 1321 -198 1323 -194
rect 1410 -189 1412 -185
rect 1430 -198 1432 -194
rect 1440 -196 1442 -191
rect 1450 -193 1452 -188
rect 1460 -193 1462 -188
rect 1498 -180 1500 -171
rect 1520 -180 1522 -171
rect 1531 -174 1533 -171
rect 1538 -174 1540 -171
rect 1558 -174 1560 -171
rect 1568 -174 1570 -171
rect 1578 -166 1580 -164
rect 1582 -166 1584 -164
rect 1578 -168 1584 -166
rect 1578 -181 1580 -168
rect 1588 -172 1590 -159
rect 1605 -160 1611 -158
rect 1605 -162 1607 -160
rect 1609 -162 1611 -160
rect 1605 -164 1611 -162
rect 1584 -174 1590 -172
rect 1609 -174 1611 -164
rect 1616 -165 1618 -155
rect 1677 -143 1679 -139
rect 1657 -157 1659 -154
rect 1653 -159 1659 -157
rect 1653 -161 1655 -159
rect 1657 -161 1659 -159
rect 1629 -165 1631 -162
rect 1653 -163 1659 -161
rect 1615 -167 1621 -165
rect 1615 -169 1617 -167
rect 1619 -169 1621 -167
rect 1615 -171 1621 -169
rect 1625 -167 1631 -165
rect 1625 -169 1627 -167
rect 1629 -169 1631 -167
rect 1625 -171 1631 -169
rect 1619 -174 1621 -171
rect 1629 -174 1631 -171
rect 1584 -176 1586 -174
rect 1588 -176 1590 -174
rect 1584 -178 1590 -176
rect 1588 -181 1590 -178
rect 1558 -193 1560 -188
rect 1568 -193 1570 -188
rect 1480 -198 1482 -194
rect 1487 -198 1489 -194
rect 1498 -198 1500 -194
rect 1520 -198 1522 -194
rect 1531 -198 1533 -194
rect 1538 -198 1540 -194
rect 1578 -196 1580 -191
rect 1609 -185 1611 -180
rect 1619 -185 1621 -180
rect 1657 -176 1659 -163
rect 1667 -165 1669 -154
rect 1720 -137 1722 -132
rect 1727 -137 1729 -132
rect 1745 -134 1747 -130
rect 1755 -134 1757 -130
rect 1765 -134 1767 -130
rect 1787 -134 1789 -130
rect 1797 -134 1799 -130
rect 1807 -134 1809 -130
rect 1710 -146 1712 -141
rect 1677 -165 1679 -161
rect 1663 -167 1669 -165
rect 1663 -169 1665 -167
rect 1667 -169 1669 -167
rect 1663 -171 1669 -169
rect 1673 -167 1679 -165
rect 1673 -169 1675 -167
rect 1677 -169 1679 -167
rect 1673 -171 1679 -169
rect 1664 -176 1666 -171
rect 1677 -176 1679 -171
rect 1697 -172 1699 -159
rect 1710 -162 1712 -159
rect 1825 -137 1827 -132
rect 1832 -137 1834 -132
rect 1855 -134 1857 -130
rect 1876 -134 1878 -130
rect 1883 -134 1885 -130
rect 1842 -146 1844 -141
rect 1927 -134 1929 -130
rect 1896 -144 1898 -139
rect 1876 -158 1878 -155
rect 1842 -162 1844 -159
rect 1703 -164 1712 -162
rect 1703 -166 1705 -164
rect 1707 -166 1709 -164
rect 1720 -165 1722 -162
rect 1727 -165 1729 -162
rect 1745 -165 1747 -162
rect 1755 -165 1757 -162
rect 1765 -165 1767 -162
rect 1787 -165 1789 -162
rect 1797 -165 1799 -162
rect 1807 -165 1809 -162
rect 1825 -165 1827 -162
rect 1832 -165 1834 -162
rect 1842 -164 1851 -162
rect 1703 -168 1709 -166
rect 1697 -174 1703 -172
rect 1697 -176 1699 -174
rect 1701 -176 1703 -174
rect 1629 -188 1631 -183
rect 1697 -178 1703 -176
rect 1697 -181 1699 -178
rect 1707 -181 1709 -168
rect 1717 -167 1723 -165
rect 1717 -169 1719 -167
rect 1721 -169 1723 -167
rect 1717 -171 1723 -169
rect 1727 -167 1749 -165
rect 1727 -169 1738 -167
rect 1740 -169 1745 -167
rect 1747 -169 1749 -167
rect 1727 -171 1749 -169
rect 1753 -167 1759 -165
rect 1753 -169 1755 -167
rect 1757 -169 1759 -167
rect 1753 -171 1759 -169
rect 1763 -167 1769 -165
rect 1763 -169 1765 -167
rect 1767 -169 1769 -167
rect 1763 -171 1769 -169
rect 1785 -167 1791 -165
rect 1785 -169 1787 -167
rect 1789 -169 1791 -167
rect 1785 -171 1791 -169
rect 1795 -167 1801 -165
rect 1795 -169 1797 -167
rect 1799 -169 1801 -167
rect 1795 -171 1801 -169
rect 1805 -167 1827 -165
rect 1805 -169 1807 -167
rect 1809 -169 1814 -167
rect 1816 -169 1827 -167
rect 1805 -171 1827 -169
rect 1831 -167 1837 -165
rect 1831 -169 1833 -167
rect 1835 -169 1837 -167
rect 1831 -171 1837 -169
rect 1717 -174 1719 -171
rect 1727 -174 1729 -171
rect 1747 -174 1749 -171
rect 1754 -174 1756 -171
rect 1657 -192 1659 -187
rect 1664 -192 1666 -187
rect 1588 -198 1590 -194
rect 1677 -189 1679 -185
rect 1697 -198 1699 -194
rect 1707 -196 1709 -191
rect 1717 -193 1719 -188
rect 1727 -193 1729 -188
rect 1765 -180 1767 -171
rect 1787 -180 1789 -171
rect 1798 -174 1800 -171
rect 1805 -174 1807 -171
rect 1825 -174 1827 -171
rect 1835 -174 1837 -171
rect 1845 -166 1847 -164
rect 1849 -166 1851 -164
rect 1845 -168 1851 -166
rect 1845 -181 1847 -168
rect 1855 -172 1857 -159
rect 1872 -160 1878 -158
rect 1872 -162 1874 -160
rect 1876 -162 1878 -160
rect 1872 -164 1878 -162
rect 1851 -174 1857 -172
rect 1876 -174 1878 -164
rect 1883 -165 1885 -155
rect 1912 -159 1918 -157
rect 1912 -161 1914 -159
rect 1916 -161 1918 -159
rect 1963 -134 1965 -130
rect 1983 -134 1985 -130
rect 1943 -143 1945 -139
rect 1953 -143 1955 -139
rect 2006 -137 2008 -132
rect 2013 -137 2015 -132
rect 2031 -134 2033 -130
rect 2041 -134 2043 -130
rect 2051 -134 2053 -130
rect 2073 -134 2075 -130
rect 2083 -134 2085 -130
rect 2093 -134 2095 -130
rect 1996 -146 1998 -141
rect 1896 -165 1898 -162
rect 1912 -163 1918 -161
rect 1882 -167 1888 -165
rect 1882 -169 1884 -167
rect 1886 -169 1888 -167
rect 1882 -171 1888 -169
rect 1892 -167 1898 -165
rect 1916 -164 1918 -163
rect 1927 -164 1929 -161
rect 1943 -164 1945 -161
rect 1916 -166 1929 -164
rect 1935 -166 1945 -164
rect 1953 -165 1955 -161
rect 1963 -164 1965 -161
rect 1892 -169 1894 -167
rect 1896 -169 1898 -167
rect 1892 -171 1898 -169
rect 1886 -174 1888 -171
rect 1896 -174 1898 -171
rect 1919 -174 1921 -166
rect 1935 -170 1937 -166
rect 1928 -172 1937 -170
rect 1949 -167 1955 -165
rect 1949 -169 1951 -167
rect 1953 -169 1955 -167
rect 1949 -171 1955 -169
rect 1959 -166 1965 -164
rect 1959 -168 1961 -166
rect 1963 -168 1965 -166
rect 1959 -170 1965 -168
rect 1928 -174 1930 -172
rect 1932 -174 1937 -172
rect 1851 -176 1853 -174
rect 1855 -176 1857 -174
rect 1851 -178 1857 -176
rect 1855 -181 1857 -178
rect 1825 -193 1827 -188
rect 1835 -193 1837 -188
rect 1747 -198 1749 -194
rect 1754 -198 1756 -194
rect 1765 -198 1767 -194
rect 1787 -198 1789 -194
rect 1798 -198 1800 -194
rect 1805 -198 1807 -194
rect 1845 -196 1847 -191
rect 1876 -185 1878 -180
rect 1886 -185 1888 -180
rect 1928 -176 1937 -174
rect 1953 -174 1955 -171
rect 1935 -179 1937 -176
rect 1945 -179 1947 -175
rect 1953 -176 1957 -174
rect 1955 -179 1957 -176
rect 1962 -179 1964 -170
rect 1983 -172 1985 -159
rect 1996 -162 1998 -159
rect 2111 -137 2113 -132
rect 2118 -137 2120 -132
rect 2141 -134 2143 -130
rect 2162 -134 2164 -130
rect 2169 -134 2171 -130
rect 2128 -146 2130 -141
rect 2216 -134 2218 -130
rect 2223 -134 2225 -130
rect 2233 -134 2235 -130
rect 2240 -134 2242 -130
rect 2250 -134 2252 -130
rect 2284 -134 2286 -130
rect 2291 -134 2293 -130
rect 2301 -134 2303 -130
rect 2308 -134 2310 -130
rect 2318 -134 2320 -130
rect 2182 -144 2184 -139
rect 2162 -158 2164 -155
rect 2128 -162 2130 -159
rect 1989 -164 1998 -162
rect 1989 -166 1991 -164
rect 1993 -166 1995 -164
rect 2006 -165 2008 -162
rect 2013 -165 2015 -162
rect 2031 -165 2033 -162
rect 2041 -165 2043 -162
rect 2051 -165 2053 -162
rect 2073 -165 2075 -162
rect 2083 -165 2085 -162
rect 2093 -165 2095 -162
rect 2111 -165 2113 -162
rect 2118 -165 2120 -162
rect 2128 -164 2137 -162
rect 1989 -168 1995 -166
rect 1983 -174 1989 -172
rect 1983 -176 1985 -174
rect 1987 -176 1989 -174
rect 1983 -178 1989 -176
rect 1896 -188 1898 -183
rect 1919 -186 1921 -183
rect 1919 -188 1924 -186
rect 1855 -198 1857 -194
rect 1922 -196 1924 -188
rect 1935 -192 1937 -188
rect 1945 -196 1947 -188
rect 1983 -181 1985 -178
rect 1993 -181 1995 -168
rect 2003 -167 2009 -165
rect 2003 -169 2005 -167
rect 2007 -169 2009 -167
rect 2003 -171 2009 -169
rect 2013 -167 2035 -165
rect 2013 -169 2024 -167
rect 2026 -169 2031 -167
rect 2033 -169 2035 -167
rect 2013 -171 2035 -169
rect 2039 -167 2045 -165
rect 2039 -169 2041 -167
rect 2043 -169 2045 -167
rect 2039 -171 2045 -169
rect 2049 -167 2055 -165
rect 2049 -169 2051 -167
rect 2053 -169 2055 -167
rect 2049 -171 2055 -169
rect 2071 -167 2077 -165
rect 2071 -169 2073 -167
rect 2075 -169 2077 -167
rect 2071 -171 2077 -169
rect 2081 -167 2087 -165
rect 2081 -169 2083 -167
rect 2085 -169 2087 -167
rect 2081 -171 2087 -169
rect 2091 -167 2113 -165
rect 2091 -169 2093 -167
rect 2095 -169 2100 -167
rect 2102 -169 2113 -167
rect 2091 -171 2113 -169
rect 2117 -167 2123 -165
rect 2117 -169 2119 -167
rect 2121 -169 2123 -167
rect 2117 -171 2123 -169
rect 2003 -174 2005 -171
rect 2013 -174 2015 -171
rect 2033 -174 2035 -171
rect 2040 -174 2042 -171
rect 1955 -196 1957 -191
rect 1962 -196 1964 -191
rect 1922 -198 1947 -196
rect 1983 -198 1985 -194
rect 1993 -196 1995 -191
rect 2003 -193 2005 -188
rect 2013 -193 2015 -188
rect 2051 -180 2053 -171
rect 2073 -180 2075 -171
rect 2084 -174 2086 -171
rect 2091 -174 2093 -171
rect 2111 -174 2113 -171
rect 2121 -174 2123 -171
rect 2131 -166 2133 -164
rect 2135 -166 2137 -164
rect 2131 -168 2137 -166
rect 2131 -181 2133 -168
rect 2141 -172 2143 -159
rect 2158 -160 2164 -158
rect 2158 -162 2160 -160
rect 2162 -162 2164 -160
rect 2158 -164 2164 -162
rect 2137 -174 2143 -172
rect 2162 -174 2164 -164
rect 2169 -165 2171 -155
rect 2199 -147 2205 -145
rect 2199 -149 2201 -147
rect 2203 -149 2205 -147
rect 2199 -151 2208 -149
rect 2206 -154 2208 -151
rect 2182 -165 2184 -162
rect 2168 -167 2174 -165
rect 2168 -169 2170 -167
rect 2172 -169 2174 -167
rect 2168 -171 2174 -169
rect 2178 -167 2184 -165
rect 2178 -169 2180 -167
rect 2182 -169 2184 -167
rect 2178 -171 2184 -169
rect 2172 -174 2174 -171
rect 2182 -174 2184 -171
rect 2137 -176 2139 -174
rect 2141 -176 2143 -174
rect 2137 -178 2143 -176
rect 2141 -181 2143 -178
rect 2111 -193 2113 -188
rect 2121 -193 2123 -188
rect 2033 -198 2035 -194
rect 2040 -198 2042 -194
rect 2051 -198 2053 -194
rect 2073 -198 2075 -194
rect 2084 -198 2086 -194
rect 2091 -198 2093 -194
rect 2131 -196 2133 -191
rect 2162 -185 2164 -180
rect 2172 -185 2174 -180
rect 2206 -180 2208 -162
rect 2216 -165 2218 -150
rect 2223 -155 2225 -150
rect 2222 -157 2228 -155
rect 2222 -159 2224 -157
rect 2226 -159 2228 -157
rect 2222 -161 2228 -159
rect 2233 -165 2235 -150
rect 2240 -160 2242 -150
rect 2267 -147 2273 -145
rect 2267 -149 2269 -147
rect 2271 -149 2273 -147
rect 2267 -151 2276 -149
rect 2212 -167 2218 -165
rect 2212 -169 2214 -167
rect 2216 -169 2218 -167
rect 2212 -171 2218 -169
rect 2216 -180 2218 -171
rect 2223 -167 2235 -165
rect 2239 -162 2245 -160
rect 2239 -164 2241 -162
rect 2243 -164 2245 -162
rect 2239 -166 2245 -164
rect 2223 -180 2225 -167
rect 2229 -173 2235 -171
rect 2229 -175 2231 -173
rect 2233 -175 2235 -173
rect 2229 -177 2235 -175
rect 2233 -180 2235 -177
rect 2240 -180 2242 -166
rect 2250 -170 2252 -152
rect 2274 -154 2276 -151
rect 2247 -172 2253 -170
rect 2247 -174 2249 -172
rect 2251 -174 2253 -172
rect 2247 -176 2253 -174
rect 2250 -179 2252 -176
rect 2182 -188 2184 -183
rect 2141 -198 2143 -194
rect 2206 -196 2208 -186
rect 2274 -180 2276 -162
rect 2284 -165 2286 -150
rect 2291 -155 2293 -150
rect 2290 -157 2296 -155
rect 2290 -159 2292 -157
rect 2294 -159 2296 -157
rect 2290 -161 2296 -159
rect 2301 -165 2303 -150
rect 2308 -160 2310 -150
rect 2280 -167 2286 -165
rect 2280 -169 2282 -167
rect 2284 -169 2286 -167
rect 2280 -171 2286 -169
rect 2284 -180 2286 -171
rect 2291 -167 2303 -165
rect 2307 -162 2313 -160
rect 2307 -164 2309 -162
rect 2311 -164 2313 -162
rect 2307 -166 2313 -164
rect 2291 -180 2293 -167
rect 2297 -173 2303 -171
rect 2297 -175 2299 -173
rect 2301 -175 2303 -173
rect 2297 -177 2303 -175
rect 2301 -180 2303 -177
rect 2308 -180 2310 -166
rect 2318 -170 2320 -152
rect 2315 -172 2321 -170
rect 2315 -174 2317 -172
rect 2319 -174 2321 -172
rect 2315 -176 2321 -174
rect 2318 -179 2320 -176
rect 2216 -192 2218 -188
rect 2223 -196 2225 -188
rect 2233 -193 2235 -188
rect 2240 -193 2242 -188
rect 2250 -193 2252 -188
rect 2206 -198 2225 -196
rect 2274 -196 2276 -186
rect 2284 -192 2286 -188
rect 2291 -196 2293 -188
rect 2301 -193 2303 -188
rect 2308 -193 2310 -188
rect 2318 -193 2320 -188
rect 2274 -198 2293 -196
rect 15 -213 17 -208
rect 22 -213 24 -208
rect 35 -215 37 -211
rect 55 -213 57 -208
rect 62 -213 64 -208
rect 95 -206 97 -202
rect 75 -215 77 -211
rect 105 -209 107 -204
rect 145 -206 147 -202
rect 152 -206 154 -202
rect 163 -206 165 -202
rect 185 -206 187 -202
rect 196 -206 198 -202
rect 203 -206 205 -202
rect 115 -212 117 -207
rect 125 -212 127 -207
rect 95 -222 97 -219
rect 95 -224 101 -222
rect 15 -237 17 -224
rect 22 -229 24 -224
rect 35 -229 37 -224
rect 21 -231 27 -229
rect 21 -233 23 -231
rect 25 -233 27 -231
rect 21 -235 27 -233
rect 31 -231 37 -229
rect 31 -233 33 -231
rect 35 -233 37 -231
rect 31 -235 37 -233
rect 11 -239 17 -237
rect 11 -241 13 -239
rect 15 -241 17 -239
rect 11 -243 17 -241
rect 15 -246 17 -243
rect 25 -246 27 -235
rect 35 -239 37 -235
rect 55 -237 57 -224
rect 62 -229 64 -224
rect 75 -229 77 -224
rect 61 -231 67 -229
rect 61 -233 63 -231
rect 65 -233 67 -231
rect 61 -235 67 -233
rect 71 -231 77 -229
rect 71 -233 73 -231
rect 75 -233 77 -231
rect 71 -235 77 -233
rect 51 -239 57 -237
rect 51 -241 53 -239
rect 55 -241 57 -239
rect 51 -243 57 -241
rect 55 -246 57 -243
rect 65 -246 67 -235
rect 75 -239 77 -235
rect 95 -226 97 -224
rect 99 -226 101 -224
rect 95 -228 101 -226
rect 15 -264 17 -259
rect 25 -264 27 -259
rect 35 -261 37 -257
rect 95 -241 97 -228
rect 105 -232 107 -219
rect 101 -234 107 -232
rect 101 -236 103 -234
rect 105 -236 107 -234
rect 115 -229 117 -226
rect 125 -229 127 -226
rect 145 -229 147 -226
rect 152 -229 154 -226
rect 163 -229 165 -220
rect 185 -229 187 -220
rect 223 -212 225 -207
rect 233 -212 235 -207
rect 243 -209 245 -204
rect 253 -206 255 -202
rect 196 -229 198 -226
rect 203 -229 205 -226
rect 223 -229 225 -226
rect 233 -229 235 -226
rect 115 -231 121 -229
rect 115 -233 117 -231
rect 119 -233 121 -231
rect 115 -235 121 -233
rect 125 -231 147 -229
rect 125 -233 136 -231
rect 138 -233 143 -231
rect 145 -233 147 -231
rect 125 -235 147 -233
rect 151 -231 157 -229
rect 151 -233 153 -231
rect 155 -233 157 -231
rect 151 -235 157 -233
rect 161 -231 167 -229
rect 161 -233 163 -231
rect 165 -233 167 -231
rect 161 -235 167 -233
rect 183 -231 189 -229
rect 183 -233 185 -231
rect 187 -233 189 -231
rect 183 -235 189 -233
rect 193 -231 199 -229
rect 193 -233 195 -231
rect 197 -233 199 -231
rect 193 -235 199 -233
rect 203 -231 225 -229
rect 203 -233 205 -231
rect 207 -233 212 -231
rect 214 -233 225 -231
rect 203 -235 225 -233
rect 229 -231 235 -229
rect 229 -233 231 -231
rect 233 -233 235 -231
rect 229 -235 235 -233
rect 243 -232 245 -219
rect 253 -222 255 -219
rect 249 -224 255 -222
rect 249 -226 251 -224
rect 253 -226 255 -224
rect 274 -220 276 -215
rect 284 -220 286 -215
rect 294 -217 296 -212
rect 322 -213 324 -208
rect 329 -213 331 -208
rect 362 -206 364 -202
rect 342 -215 344 -211
rect 372 -209 374 -204
rect 412 -206 414 -202
rect 419 -206 421 -202
rect 430 -206 432 -202
rect 452 -206 454 -202
rect 463 -206 465 -202
rect 470 -206 472 -202
rect 382 -212 384 -207
rect 392 -212 394 -207
rect 362 -222 364 -219
rect 362 -224 368 -222
rect 249 -228 255 -226
rect 243 -234 249 -232
rect 101 -238 110 -236
rect 118 -238 120 -235
rect 125 -238 127 -235
rect 143 -238 145 -235
rect 153 -238 155 -235
rect 163 -238 165 -235
rect 185 -238 187 -235
rect 195 -238 197 -235
rect 205 -238 207 -235
rect 223 -238 225 -235
rect 230 -238 232 -235
rect 243 -236 245 -234
rect 247 -236 249 -234
rect 240 -238 249 -236
rect 108 -241 110 -238
rect 55 -264 57 -259
rect 65 -264 67 -259
rect 75 -261 77 -257
rect 108 -259 110 -254
rect 95 -270 97 -266
rect 118 -268 120 -263
rect 125 -268 127 -263
rect 240 -241 242 -238
rect 253 -241 255 -228
rect 274 -236 276 -226
rect 284 -229 286 -226
rect 294 -229 296 -226
rect 280 -231 286 -229
rect 280 -233 282 -231
rect 284 -233 286 -231
rect 280 -235 286 -233
rect 290 -231 296 -229
rect 290 -233 292 -231
rect 294 -233 296 -231
rect 290 -235 296 -233
rect 270 -238 276 -236
rect 270 -240 272 -238
rect 274 -240 276 -238
rect 240 -259 242 -254
rect 143 -270 145 -266
rect 153 -270 155 -266
rect 163 -270 165 -266
rect 185 -270 187 -266
rect 195 -270 197 -266
rect 205 -270 207 -266
rect 223 -268 225 -263
rect 230 -268 232 -263
rect 270 -242 276 -240
rect 274 -245 276 -242
rect 281 -245 283 -235
rect 294 -238 296 -235
rect 322 -237 324 -224
rect 329 -229 331 -224
rect 342 -229 344 -224
rect 328 -231 334 -229
rect 328 -233 330 -231
rect 332 -233 334 -231
rect 328 -235 334 -233
rect 338 -231 344 -229
rect 338 -233 340 -231
rect 342 -233 344 -231
rect 338 -235 344 -233
rect 318 -239 324 -237
rect 318 -241 320 -239
rect 322 -241 324 -239
rect 318 -243 324 -241
rect 322 -246 324 -243
rect 332 -246 334 -235
rect 342 -239 344 -235
rect 362 -226 364 -224
rect 366 -226 368 -224
rect 362 -228 368 -226
rect 294 -261 296 -256
rect 362 -241 364 -228
rect 372 -232 374 -219
rect 368 -234 374 -232
rect 368 -236 370 -234
rect 372 -236 374 -234
rect 382 -229 384 -226
rect 392 -229 394 -226
rect 412 -229 414 -226
rect 419 -229 421 -226
rect 430 -229 432 -220
rect 452 -229 454 -220
rect 490 -212 492 -207
rect 500 -212 502 -207
rect 510 -209 512 -204
rect 520 -206 522 -202
rect 463 -229 465 -226
rect 470 -229 472 -226
rect 490 -229 492 -226
rect 500 -229 502 -226
rect 382 -231 388 -229
rect 382 -233 384 -231
rect 386 -233 388 -231
rect 382 -235 388 -233
rect 392 -231 414 -229
rect 392 -233 403 -231
rect 405 -233 410 -231
rect 412 -233 414 -231
rect 392 -235 414 -233
rect 418 -231 424 -229
rect 418 -233 420 -231
rect 422 -233 424 -231
rect 418 -235 424 -233
rect 428 -231 434 -229
rect 428 -233 430 -231
rect 432 -233 434 -231
rect 428 -235 434 -233
rect 450 -231 456 -229
rect 450 -233 452 -231
rect 454 -233 456 -231
rect 450 -235 456 -233
rect 460 -231 466 -229
rect 460 -233 462 -231
rect 464 -233 466 -231
rect 460 -235 466 -233
rect 470 -231 492 -229
rect 470 -233 472 -231
rect 474 -233 479 -231
rect 481 -233 492 -231
rect 470 -235 492 -233
rect 496 -231 502 -229
rect 496 -233 498 -231
rect 500 -233 502 -231
rect 496 -235 502 -233
rect 510 -232 512 -219
rect 520 -222 522 -219
rect 516 -224 522 -222
rect 516 -226 518 -224
rect 520 -226 522 -224
rect 541 -220 543 -215
rect 551 -220 553 -215
rect 561 -217 563 -212
rect 589 -213 591 -208
rect 596 -213 598 -208
rect 629 -206 631 -202
rect 609 -215 611 -211
rect 639 -209 641 -204
rect 679 -206 681 -202
rect 686 -206 688 -202
rect 697 -206 699 -202
rect 719 -206 721 -202
rect 730 -206 732 -202
rect 737 -206 739 -202
rect 649 -212 651 -207
rect 659 -212 661 -207
rect 629 -222 631 -219
rect 629 -224 635 -222
rect 516 -228 522 -226
rect 510 -234 516 -232
rect 368 -238 377 -236
rect 385 -238 387 -235
rect 392 -238 394 -235
rect 410 -238 412 -235
rect 420 -238 422 -235
rect 430 -238 432 -235
rect 452 -238 454 -235
rect 462 -238 464 -235
rect 472 -238 474 -235
rect 490 -238 492 -235
rect 497 -238 499 -235
rect 510 -236 512 -234
rect 514 -236 516 -234
rect 507 -238 516 -236
rect 375 -241 377 -238
rect 322 -264 324 -259
rect 332 -264 334 -259
rect 342 -261 344 -257
rect 253 -270 255 -266
rect 274 -270 276 -266
rect 281 -270 283 -266
rect 375 -259 377 -254
rect 362 -270 364 -266
rect 385 -268 387 -263
rect 392 -268 394 -263
rect 507 -241 509 -238
rect 520 -241 522 -228
rect 541 -236 543 -226
rect 551 -229 553 -226
rect 561 -229 563 -226
rect 547 -231 553 -229
rect 547 -233 549 -231
rect 551 -233 553 -231
rect 547 -235 553 -233
rect 557 -231 563 -229
rect 557 -233 559 -231
rect 561 -233 563 -231
rect 557 -235 563 -233
rect 537 -238 543 -236
rect 537 -240 539 -238
rect 541 -240 543 -238
rect 507 -259 509 -254
rect 410 -270 412 -266
rect 420 -270 422 -266
rect 430 -270 432 -266
rect 452 -270 454 -266
rect 462 -270 464 -266
rect 472 -270 474 -266
rect 490 -268 492 -263
rect 497 -268 499 -263
rect 537 -242 543 -240
rect 541 -245 543 -242
rect 548 -245 550 -235
rect 561 -238 563 -235
rect 589 -237 591 -224
rect 596 -229 598 -224
rect 609 -229 611 -224
rect 595 -231 601 -229
rect 595 -233 597 -231
rect 599 -233 601 -231
rect 595 -235 601 -233
rect 605 -231 611 -229
rect 605 -233 607 -231
rect 609 -233 611 -231
rect 605 -235 611 -233
rect 585 -239 591 -237
rect 585 -241 587 -239
rect 589 -241 591 -239
rect 585 -243 591 -241
rect 589 -246 591 -243
rect 599 -246 601 -235
rect 609 -239 611 -235
rect 629 -226 631 -224
rect 633 -226 635 -224
rect 629 -228 635 -226
rect 561 -261 563 -256
rect 629 -241 631 -228
rect 639 -232 641 -219
rect 635 -234 641 -232
rect 635 -236 637 -234
rect 639 -236 641 -234
rect 649 -229 651 -226
rect 659 -229 661 -226
rect 679 -229 681 -226
rect 686 -229 688 -226
rect 697 -229 699 -220
rect 719 -229 721 -220
rect 757 -212 759 -207
rect 767 -212 769 -207
rect 777 -209 779 -204
rect 787 -206 789 -202
rect 730 -229 732 -226
rect 737 -229 739 -226
rect 757 -229 759 -226
rect 767 -229 769 -226
rect 649 -231 655 -229
rect 649 -233 651 -231
rect 653 -233 655 -231
rect 649 -235 655 -233
rect 659 -231 681 -229
rect 659 -233 670 -231
rect 672 -233 677 -231
rect 679 -233 681 -231
rect 659 -235 681 -233
rect 685 -231 691 -229
rect 685 -233 687 -231
rect 689 -233 691 -231
rect 685 -235 691 -233
rect 695 -231 701 -229
rect 695 -233 697 -231
rect 699 -233 701 -231
rect 695 -235 701 -233
rect 717 -231 723 -229
rect 717 -233 719 -231
rect 721 -233 723 -231
rect 717 -235 723 -233
rect 727 -231 733 -229
rect 727 -233 729 -231
rect 731 -233 733 -231
rect 727 -235 733 -233
rect 737 -231 759 -229
rect 737 -233 739 -231
rect 741 -233 746 -231
rect 748 -233 759 -231
rect 737 -235 759 -233
rect 763 -231 769 -229
rect 763 -233 765 -231
rect 767 -233 769 -231
rect 763 -235 769 -233
rect 777 -232 779 -219
rect 787 -222 789 -219
rect 783 -224 789 -222
rect 783 -226 785 -224
rect 787 -226 789 -224
rect 808 -220 810 -215
rect 818 -220 820 -215
rect 828 -217 830 -212
rect 856 -213 858 -208
rect 863 -213 865 -208
rect 896 -206 898 -202
rect 876 -215 878 -211
rect 906 -209 908 -204
rect 946 -206 948 -202
rect 953 -206 955 -202
rect 964 -206 966 -202
rect 986 -206 988 -202
rect 997 -206 999 -202
rect 1004 -206 1006 -202
rect 916 -212 918 -207
rect 926 -212 928 -207
rect 896 -222 898 -219
rect 896 -224 902 -222
rect 783 -228 789 -226
rect 777 -234 783 -232
rect 635 -238 644 -236
rect 652 -238 654 -235
rect 659 -238 661 -235
rect 677 -238 679 -235
rect 687 -238 689 -235
rect 697 -238 699 -235
rect 719 -238 721 -235
rect 729 -238 731 -235
rect 739 -238 741 -235
rect 757 -238 759 -235
rect 764 -238 766 -235
rect 777 -236 779 -234
rect 781 -236 783 -234
rect 774 -238 783 -236
rect 642 -241 644 -238
rect 589 -264 591 -259
rect 599 -264 601 -259
rect 609 -261 611 -257
rect 520 -270 522 -266
rect 541 -270 543 -266
rect 548 -270 550 -266
rect 642 -259 644 -254
rect 629 -270 631 -266
rect 652 -268 654 -263
rect 659 -268 661 -263
rect 774 -241 776 -238
rect 787 -241 789 -228
rect 808 -236 810 -226
rect 818 -229 820 -226
rect 828 -229 830 -226
rect 814 -231 820 -229
rect 814 -233 816 -231
rect 818 -233 820 -231
rect 814 -235 820 -233
rect 824 -231 830 -229
rect 824 -233 826 -231
rect 828 -233 830 -231
rect 824 -235 830 -233
rect 804 -238 810 -236
rect 804 -240 806 -238
rect 808 -240 810 -238
rect 774 -259 776 -254
rect 677 -270 679 -266
rect 687 -270 689 -266
rect 697 -270 699 -266
rect 719 -270 721 -266
rect 729 -270 731 -266
rect 739 -270 741 -266
rect 757 -268 759 -263
rect 764 -268 766 -263
rect 804 -242 810 -240
rect 808 -245 810 -242
rect 815 -245 817 -235
rect 828 -238 830 -235
rect 856 -237 858 -224
rect 863 -229 865 -224
rect 876 -229 878 -224
rect 862 -231 868 -229
rect 862 -233 864 -231
rect 866 -233 868 -231
rect 862 -235 868 -233
rect 872 -231 878 -229
rect 872 -233 874 -231
rect 876 -233 878 -231
rect 872 -235 878 -233
rect 852 -239 858 -237
rect 852 -241 854 -239
rect 856 -241 858 -239
rect 852 -243 858 -241
rect 856 -246 858 -243
rect 866 -246 868 -235
rect 876 -239 878 -235
rect 896 -226 898 -224
rect 900 -226 902 -224
rect 896 -228 902 -226
rect 828 -261 830 -256
rect 896 -241 898 -228
rect 906 -232 908 -219
rect 902 -234 908 -232
rect 902 -236 904 -234
rect 906 -236 908 -234
rect 916 -229 918 -226
rect 926 -229 928 -226
rect 946 -229 948 -226
rect 953 -229 955 -226
rect 964 -229 966 -220
rect 986 -229 988 -220
rect 1024 -212 1026 -207
rect 1034 -212 1036 -207
rect 1044 -209 1046 -204
rect 1054 -206 1056 -202
rect 997 -229 999 -226
rect 1004 -229 1006 -226
rect 1024 -229 1026 -226
rect 1034 -229 1036 -226
rect 916 -231 922 -229
rect 916 -233 918 -231
rect 920 -233 922 -231
rect 916 -235 922 -233
rect 926 -231 948 -229
rect 926 -233 937 -231
rect 939 -233 944 -231
rect 946 -233 948 -231
rect 926 -235 948 -233
rect 952 -231 958 -229
rect 952 -233 954 -231
rect 956 -233 958 -231
rect 952 -235 958 -233
rect 962 -231 968 -229
rect 962 -233 964 -231
rect 966 -233 968 -231
rect 962 -235 968 -233
rect 984 -231 990 -229
rect 984 -233 986 -231
rect 988 -233 990 -231
rect 984 -235 990 -233
rect 994 -231 1000 -229
rect 994 -233 996 -231
rect 998 -233 1000 -231
rect 994 -235 1000 -233
rect 1004 -231 1026 -229
rect 1004 -233 1006 -231
rect 1008 -233 1013 -231
rect 1015 -233 1026 -231
rect 1004 -235 1026 -233
rect 1030 -231 1036 -229
rect 1030 -233 1032 -231
rect 1034 -233 1036 -231
rect 1030 -235 1036 -233
rect 1044 -232 1046 -219
rect 1054 -222 1056 -219
rect 1050 -224 1056 -222
rect 1050 -226 1052 -224
rect 1054 -226 1056 -224
rect 1075 -220 1077 -215
rect 1085 -220 1087 -215
rect 1095 -217 1097 -212
rect 1123 -213 1125 -208
rect 1130 -213 1132 -208
rect 1163 -206 1165 -202
rect 1143 -215 1145 -211
rect 1173 -209 1175 -204
rect 1213 -206 1215 -202
rect 1220 -206 1222 -202
rect 1231 -206 1233 -202
rect 1253 -206 1255 -202
rect 1264 -206 1266 -202
rect 1271 -206 1273 -202
rect 1183 -212 1185 -207
rect 1193 -212 1195 -207
rect 1163 -222 1165 -219
rect 1163 -224 1169 -222
rect 1050 -228 1056 -226
rect 1044 -234 1050 -232
rect 902 -238 911 -236
rect 919 -238 921 -235
rect 926 -238 928 -235
rect 944 -238 946 -235
rect 954 -238 956 -235
rect 964 -238 966 -235
rect 986 -238 988 -235
rect 996 -238 998 -235
rect 1006 -238 1008 -235
rect 1024 -238 1026 -235
rect 1031 -238 1033 -235
rect 1044 -236 1046 -234
rect 1048 -236 1050 -234
rect 1041 -238 1050 -236
rect 909 -241 911 -238
rect 856 -264 858 -259
rect 866 -264 868 -259
rect 876 -261 878 -257
rect 787 -270 789 -266
rect 808 -270 810 -266
rect 815 -270 817 -266
rect 909 -259 911 -254
rect 896 -270 898 -266
rect 919 -268 921 -263
rect 926 -268 928 -263
rect 1041 -241 1043 -238
rect 1054 -241 1056 -228
rect 1075 -236 1077 -226
rect 1085 -229 1087 -226
rect 1095 -229 1097 -226
rect 1081 -231 1087 -229
rect 1081 -233 1083 -231
rect 1085 -233 1087 -231
rect 1081 -235 1087 -233
rect 1091 -231 1097 -229
rect 1091 -233 1093 -231
rect 1095 -233 1097 -231
rect 1091 -235 1097 -233
rect 1071 -238 1077 -236
rect 1071 -240 1073 -238
rect 1075 -240 1077 -238
rect 1041 -259 1043 -254
rect 944 -270 946 -266
rect 954 -270 956 -266
rect 964 -270 966 -266
rect 986 -270 988 -266
rect 996 -270 998 -266
rect 1006 -270 1008 -266
rect 1024 -268 1026 -263
rect 1031 -268 1033 -263
rect 1071 -242 1077 -240
rect 1075 -245 1077 -242
rect 1082 -245 1084 -235
rect 1095 -238 1097 -235
rect 1123 -237 1125 -224
rect 1130 -229 1132 -224
rect 1143 -229 1145 -224
rect 1129 -231 1135 -229
rect 1129 -233 1131 -231
rect 1133 -233 1135 -231
rect 1129 -235 1135 -233
rect 1139 -231 1145 -229
rect 1139 -233 1141 -231
rect 1143 -233 1145 -231
rect 1139 -235 1145 -233
rect 1119 -239 1125 -237
rect 1119 -241 1121 -239
rect 1123 -241 1125 -239
rect 1119 -243 1125 -241
rect 1123 -246 1125 -243
rect 1133 -246 1135 -235
rect 1143 -239 1145 -235
rect 1163 -226 1165 -224
rect 1167 -226 1169 -224
rect 1163 -228 1169 -226
rect 1095 -261 1097 -256
rect 1163 -241 1165 -228
rect 1173 -232 1175 -219
rect 1169 -234 1175 -232
rect 1169 -236 1171 -234
rect 1173 -236 1175 -234
rect 1183 -229 1185 -226
rect 1193 -229 1195 -226
rect 1213 -229 1215 -226
rect 1220 -229 1222 -226
rect 1231 -229 1233 -220
rect 1253 -229 1255 -220
rect 1291 -212 1293 -207
rect 1301 -212 1303 -207
rect 1311 -209 1313 -204
rect 1321 -206 1323 -202
rect 1264 -229 1266 -226
rect 1271 -229 1273 -226
rect 1291 -229 1293 -226
rect 1301 -229 1303 -226
rect 1183 -231 1189 -229
rect 1183 -233 1185 -231
rect 1187 -233 1189 -231
rect 1183 -235 1189 -233
rect 1193 -231 1215 -229
rect 1193 -233 1204 -231
rect 1206 -233 1211 -231
rect 1213 -233 1215 -231
rect 1193 -235 1215 -233
rect 1219 -231 1225 -229
rect 1219 -233 1221 -231
rect 1223 -233 1225 -231
rect 1219 -235 1225 -233
rect 1229 -231 1235 -229
rect 1229 -233 1231 -231
rect 1233 -233 1235 -231
rect 1229 -235 1235 -233
rect 1251 -231 1257 -229
rect 1251 -233 1253 -231
rect 1255 -233 1257 -231
rect 1251 -235 1257 -233
rect 1261 -231 1267 -229
rect 1261 -233 1263 -231
rect 1265 -233 1267 -231
rect 1261 -235 1267 -233
rect 1271 -231 1293 -229
rect 1271 -233 1273 -231
rect 1275 -233 1280 -231
rect 1282 -233 1293 -231
rect 1271 -235 1293 -233
rect 1297 -231 1303 -229
rect 1297 -233 1299 -231
rect 1301 -233 1303 -231
rect 1297 -235 1303 -233
rect 1311 -232 1313 -219
rect 1321 -222 1323 -219
rect 1317 -224 1323 -222
rect 1317 -226 1319 -224
rect 1321 -226 1323 -224
rect 1342 -220 1344 -215
rect 1352 -220 1354 -215
rect 1362 -217 1364 -212
rect 1390 -213 1392 -208
rect 1397 -213 1399 -208
rect 1430 -206 1432 -202
rect 1410 -215 1412 -211
rect 1440 -209 1442 -204
rect 1480 -206 1482 -202
rect 1487 -206 1489 -202
rect 1498 -206 1500 -202
rect 1520 -206 1522 -202
rect 1531 -206 1533 -202
rect 1538 -206 1540 -202
rect 1450 -212 1452 -207
rect 1460 -212 1462 -207
rect 1430 -222 1432 -219
rect 1430 -224 1436 -222
rect 1317 -228 1323 -226
rect 1311 -234 1317 -232
rect 1169 -238 1178 -236
rect 1186 -238 1188 -235
rect 1193 -238 1195 -235
rect 1211 -238 1213 -235
rect 1221 -238 1223 -235
rect 1231 -238 1233 -235
rect 1253 -238 1255 -235
rect 1263 -238 1265 -235
rect 1273 -238 1275 -235
rect 1291 -238 1293 -235
rect 1298 -238 1300 -235
rect 1311 -236 1313 -234
rect 1315 -236 1317 -234
rect 1308 -238 1317 -236
rect 1176 -241 1178 -238
rect 1123 -264 1125 -259
rect 1133 -264 1135 -259
rect 1143 -261 1145 -257
rect 1054 -270 1056 -266
rect 1075 -270 1077 -266
rect 1082 -270 1084 -266
rect 1176 -259 1178 -254
rect 1163 -270 1165 -266
rect 1186 -268 1188 -263
rect 1193 -268 1195 -263
rect 1308 -241 1310 -238
rect 1321 -241 1323 -228
rect 1342 -236 1344 -226
rect 1352 -229 1354 -226
rect 1362 -229 1364 -226
rect 1348 -231 1354 -229
rect 1348 -233 1350 -231
rect 1352 -233 1354 -231
rect 1348 -235 1354 -233
rect 1358 -231 1364 -229
rect 1358 -233 1360 -231
rect 1362 -233 1364 -231
rect 1358 -235 1364 -233
rect 1338 -238 1344 -236
rect 1338 -240 1340 -238
rect 1342 -240 1344 -238
rect 1308 -259 1310 -254
rect 1211 -270 1213 -266
rect 1221 -270 1223 -266
rect 1231 -270 1233 -266
rect 1253 -270 1255 -266
rect 1263 -270 1265 -266
rect 1273 -270 1275 -266
rect 1291 -268 1293 -263
rect 1298 -268 1300 -263
rect 1338 -242 1344 -240
rect 1342 -245 1344 -242
rect 1349 -245 1351 -235
rect 1362 -238 1364 -235
rect 1390 -237 1392 -224
rect 1397 -229 1399 -224
rect 1410 -229 1412 -224
rect 1396 -231 1402 -229
rect 1396 -233 1398 -231
rect 1400 -233 1402 -231
rect 1396 -235 1402 -233
rect 1406 -231 1412 -229
rect 1406 -233 1408 -231
rect 1410 -233 1412 -231
rect 1406 -235 1412 -233
rect 1386 -239 1392 -237
rect 1386 -241 1388 -239
rect 1390 -241 1392 -239
rect 1386 -243 1392 -241
rect 1390 -246 1392 -243
rect 1400 -246 1402 -235
rect 1410 -239 1412 -235
rect 1430 -226 1432 -224
rect 1434 -226 1436 -224
rect 1430 -228 1436 -226
rect 1362 -261 1364 -256
rect 1430 -241 1432 -228
rect 1440 -232 1442 -219
rect 1436 -234 1442 -232
rect 1436 -236 1438 -234
rect 1440 -236 1442 -234
rect 1450 -229 1452 -226
rect 1460 -229 1462 -226
rect 1480 -229 1482 -226
rect 1487 -229 1489 -226
rect 1498 -229 1500 -220
rect 1520 -229 1522 -220
rect 1558 -212 1560 -207
rect 1568 -212 1570 -207
rect 1578 -209 1580 -204
rect 1588 -206 1590 -202
rect 1531 -229 1533 -226
rect 1538 -229 1540 -226
rect 1558 -229 1560 -226
rect 1568 -229 1570 -226
rect 1450 -231 1456 -229
rect 1450 -233 1452 -231
rect 1454 -233 1456 -231
rect 1450 -235 1456 -233
rect 1460 -231 1482 -229
rect 1460 -233 1471 -231
rect 1473 -233 1478 -231
rect 1480 -233 1482 -231
rect 1460 -235 1482 -233
rect 1486 -231 1492 -229
rect 1486 -233 1488 -231
rect 1490 -233 1492 -231
rect 1486 -235 1492 -233
rect 1496 -231 1502 -229
rect 1496 -233 1498 -231
rect 1500 -233 1502 -231
rect 1496 -235 1502 -233
rect 1518 -231 1524 -229
rect 1518 -233 1520 -231
rect 1522 -233 1524 -231
rect 1518 -235 1524 -233
rect 1528 -231 1534 -229
rect 1528 -233 1530 -231
rect 1532 -233 1534 -231
rect 1528 -235 1534 -233
rect 1538 -231 1560 -229
rect 1538 -233 1540 -231
rect 1542 -233 1547 -231
rect 1549 -233 1560 -231
rect 1538 -235 1560 -233
rect 1564 -231 1570 -229
rect 1564 -233 1566 -231
rect 1568 -233 1570 -231
rect 1564 -235 1570 -233
rect 1578 -232 1580 -219
rect 1588 -222 1590 -219
rect 1584 -224 1590 -222
rect 1584 -226 1586 -224
rect 1588 -226 1590 -224
rect 1609 -220 1611 -215
rect 1619 -220 1621 -215
rect 1629 -217 1631 -212
rect 1657 -213 1659 -208
rect 1664 -213 1666 -208
rect 1697 -206 1699 -202
rect 1677 -215 1679 -211
rect 1707 -209 1709 -204
rect 1747 -206 1749 -202
rect 1754 -206 1756 -202
rect 1765 -206 1767 -202
rect 1787 -206 1789 -202
rect 1798 -206 1800 -202
rect 1805 -206 1807 -202
rect 1717 -212 1719 -207
rect 1727 -212 1729 -207
rect 1697 -222 1699 -219
rect 1697 -224 1703 -222
rect 1584 -228 1590 -226
rect 1578 -234 1584 -232
rect 1436 -238 1445 -236
rect 1453 -238 1455 -235
rect 1460 -238 1462 -235
rect 1478 -238 1480 -235
rect 1488 -238 1490 -235
rect 1498 -238 1500 -235
rect 1520 -238 1522 -235
rect 1530 -238 1532 -235
rect 1540 -238 1542 -235
rect 1558 -238 1560 -235
rect 1565 -238 1567 -235
rect 1578 -236 1580 -234
rect 1582 -236 1584 -234
rect 1575 -238 1584 -236
rect 1443 -241 1445 -238
rect 1390 -264 1392 -259
rect 1400 -264 1402 -259
rect 1410 -261 1412 -257
rect 1321 -270 1323 -266
rect 1342 -270 1344 -266
rect 1349 -270 1351 -266
rect 1443 -259 1445 -254
rect 1430 -270 1432 -266
rect 1453 -268 1455 -263
rect 1460 -268 1462 -263
rect 1575 -241 1577 -238
rect 1588 -241 1590 -228
rect 1609 -236 1611 -226
rect 1619 -229 1621 -226
rect 1629 -229 1631 -226
rect 1615 -231 1621 -229
rect 1615 -233 1617 -231
rect 1619 -233 1621 -231
rect 1615 -235 1621 -233
rect 1625 -231 1631 -229
rect 1625 -233 1627 -231
rect 1629 -233 1631 -231
rect 1625 -235 1631 -233
rect 1605 -238 1611 -236
rect 1605 -240 1607 -238
rect 1609 -240 1611 -238
rect 1575 -259 1577 -254
rect 1478 -270 1480 -266
rect 1488 -270 1490 -266
rect 1498 -270 1500 -266
rect 1520 -270 1522 -266
rect 1530 -270 1532 -266
rect 1540 -270 1542 -266
rect 1558 -268 1560 -263
rect 1565 -268 1567 -263
rect 1605 -242 1611 -240
rect 1609 -245 1611 -242
rect 1616 -245 1618 -235
rect 1629 -238 1631 -235
rect 1657 -237 1659 -224
rect 1664 -229 1666 -224
rect 1677 -229 1679 -224
rect 1663 -231 1669 -229
rect 1663 -233 1665 -231
rect 1667 -233 1669 -231
rect 1663 -235 1669 -233
rect 1673 -231 1679 -229
rect 1673 -233 1675 -231
rect 1677 -233 1679 -231
rect 1673 -235 1679 -233
rect 1653 -239 1659 -237
rect 1653 -241 1655 -239
rect 1657 -241 1659 -239
rect 1653 -243 1659 -241
rect 1657 -246 1659 -243
rect 1667 -246 1669 -235
rect 1677 -239 1679 -235
rect 1697 -226 1699 -224
rect 1701 -226 1703 -224
rect 1697 -228 1703 -226
rect 1629 -261 1631 -256
rect 1697 -241 1699 -228
rect 1707 -232 1709 -219
rect 1703 -234 1709 -232
rect 1703 -236 1705 -234
rect 1707 -236 1709 -234
rect 1717 -229 1719 -226
rect 1727 -229 1729 -226
rect 1747 -229 1749 -226
rect 1754 -229 1756 -226
rect 1765 -229 1767 -220
rect 1787 -229 1789 -220
rect 1825 -212 1827 -207
rect 1835 -212 1837 -207
rect 1845 -209 1847 -204
rect 1855 -206 1857 -202
rect 1922 -204 1947 -202
rect 1922 -212 1924 -204
rect 1935 -212 1937 -208
rect 1945 -212 1947 -204
rect 1955 -209 1957 -204
rect 1962 -209 1964 -204
rect 1983 -206 1985 -202
rect 1798 -229 1800 -226
rect 1805 -229 1807 -226
rect 1825 -229 1827 -226
rect 1835 -229 1837 -226
rect 1717 -231 1723 -229
rect 1717 -233 1719 -231
rect 1721 -233 1723 -231
rect 1717 -235 1723 -233
rect 1727 -231 1749 -229
rect 1727 -233 1738 -231
rect 1740 -233 1745 -231
rect 1747 -233 1749 -231
rect 1727 -235 1749 -233
rect 1753 -231 1759 -229
rect 1753 -233 1755 -231
rect 1757 -233 1759 -231
rect 1753 -235 1759 -233
rect 1763 -231 1769 -229
rect 1763 -233 1765 -231
rect 1767 -233 1769 -231
rect 1763 -235 1769 -233
rect 1785 -231 1791 -229
rect 1785 -233 1787 -231
rect 1789 -233 1791 -231
rect 1785 -235 1791 -233
rect 1795 -231 1801 -229
rect 1795 -233 1797 -231
rect 1799 -233 1801 -231
rect 1795 -235 1801 -233
rect 1805 -231 1827 -229
rect 1805 -233 1807 -231
rect 1809 -233 1814 -231
rect 1816 -233 1827 -231
rect 1805 -235 1827 -233
rect 1831 -231 1837 -229
rect 1831 -233 1833 -231
rect 1835 -233 1837 -231
rect 1831 -235 1837 -233
rect 1845 -232 1847 -219
rect 1855 -222 1857 -219
rect 1851 -224 1857 -222
rect 1851 -226 1853 -224
rect 1855 -226 1857 -224
rect 1876 -220 1878 -215
rect 1886 -220 1888 -215
rect 1896 -217 1898 -212
rect 1919 -214 1924 -212
rect 1919 -217 1921 -214
rect 1993 -209 1995 -204
rect 2033 -206 2035 -202
rect 2040 -206 2042 -202
rect 2051 -206 2053 -202
rect 2073 -206 2075 -202
rect 2084 -206 2086 -202
rect 2091 -206 2093 -202
rect 2003 -212 2005 -207
rect 2013 -212 2015 -207
rect 1935 -224 1937 -221
rect 1928 -226 1937 -224
rect 1945 -225 1947 -221
rect 1955 -224 1957 -221
rect 1851 -228 1857 -226
rect 1845 -234 1851 -232
rect 1703 -238 1712 -236
rect 1720 -238 1722 -235
rect 1727 -238 1729 -235
rect 1745 -238 1747 -235
rect 1755 -238 1757 -235
rect 1765 -238 1767 -235
rect 1787 -238 1789 -235
rect 1797 -238 1799 -235
rect 1807 -238 1809 -235
rect 1825 -238 1827 -235
rect 1832 -238 1834 -235
rect 1845 -236 1847 -234
rect 1849 -236 1851 -234
rect 1842 -238 1851 -236
rect 1710 -241 1712 -238
rect 1657 -264 1659 -259
rect 1667 -264 1669 -259
rect 1677 -261 1679 -257
rect 1588 -270 1590 -266
rect 1609 -270 1611 -266
rect 1616 -270 1618 -266
rect 1710 -259 1712 -254
rect 1697 -270 1699 -266
rect 1720 -268 1722 -263
rect 1727 -268 1729 -263
rect 1842 -241 1844 -238
rect 1855 -241 1857 -228
rect 1876 -236 1878 -226
rect 1886 -229 1888 -226
rect 1896 -229 1898 -226
rect 1882 -231 1888 -229
rect 1882 -233 1884 -231
rect 1886 -233 1888 -231
rect 1882 -235 1888 -233
rect 1892 -231 1898 -229
rect 1892 -233 1894 -231
rect 1896 -233 1898 -231
rect 1892 -235 1898 -233
rect 1919 -234 1921 -226
rect 1928 -228 1930 -226
rect 1932 -228 1937 -226
rect 1928 -230 1937 -228
rect 1953 -226 1957 -224
rect 1953 -229 1955 -226
rect 1935 -234 1937 -230
rect 1949 -231 1955 -229
rect 1962 -230 1964 -221
rect 1983 -222 1985 -219
rect 1983 -224 1989 -222
rect 1983 -226 1985 -224
rect 1987 -226 1989 -224
rect 1983 -228 1989 -226
rect 1949 -233 1951 -231
rect 1953 -233 1955 -231
rect 1872 -238 1878 -236
rect 1872 -240 1874 -238
rect 1876 -240 1878 -238
rect 1842 -259 1844 -254
rect 1745 -270 1747 -266
rect 1755 -270 1757 -266
rect 1765 -270 1767 -266
rect 1787 -270 1789 -266
rect 1797 -270 1799 -266
rect 1807 -270 1809 -266
rect 1825 -268 1827 -263
rect 1832 -268 1834 -263
rect 1872 -242 1878 -240
rect 1876 -245 1878 -242
rect 1883 -245 1885 -235
rect 1896 -238 1898 -235
rect 1916 -236 1929 -234
rect 1935 -236 1945 -234
rect 1949 -235 1955 -233
rect 1916 -237 1918 -236
rect 1912 -239 1918 -237
rect 1927 -239 1929 -236
rect 1943 -239 1945 -236
rect 1953 -239 1955 -235
rect 1959 -232 1965 -230
rect 1959 -234 1961 -232
rect 1963 -234 1965 -232
rect 1959 -236 1965 -234
rect 1963 -239 1965 -236
rect 1912 -241 1914 -239
rect 1916 -241 1918 -239
rect 1912 -243 1918 -241
rect 1896 -261 1898 -256
rect 1855 -270 1857 -266
rect 1876 -270 1878 -266
rect 1883 -270 1885 -266
rect 1943 -261 1945 -257
rect 1953 -261 1955 -257
rect 1927 -270 1929 -266
rect 1983 -241 1985 -228
rect 1993 -232 1995 -219
rect 1989 -234 1995 -232
rect 1989 -236 1991 -234
rect 1993 -236 1995 -234
rect 2003 -229 2005 -226
rect 2013 -229 2015 -226
rect 2033 -229 2035 -226
rect 2040 -229 2042 -226
rect 2051 -229 2053 -220
rect 2073 -229 2075 -220
rect 2111 -212 2113 -207
rect 2121 -212 2123 -207
rect 2131 -209 2133 -204
rect 2141 -206 2143 -202
rect 2206 -204 2225 -202
rect 2084 -229 2086 -226
rect 2091 -229 2093 -226
rect 2111 -229 2113 -226
rect 2121 -229 2123 -226
rect 2003 -231 2009 -229
rect 2003 -233 2005 -231
rect 2007 -233 2009 -231
rect 2003 -235 2009 -233
rect 2013 -231 2035 -229
rect 2013 -233 2024 -231
rect 2026 -233 2031 -231
rect 2033 -233 2035 -231
rect 2013 -235 2035 -233
rect 2039 -231 2045 -229
rect 2039 -233 2041 -231
rect 2043 -233 2045 -231
rect 2039 -235 2045 -233
rect 2049 -231 2055 -229
rect 2049 -233 2051 -231
rect 2053 -233 2055 -231
rect 2049 -235 2055 -233
rect 2071 -231 2077 -229
rect 2071 -233 2073 -231
rect 2075 -233 2077 -231
rect 2071 -235 2077 -233
rect 2081 -231 2087 -229
rect 2081 -233 2083 -231
rect 2085 -233 2087 -231
rect 2081 -235 2087 -233
rect 2091 -231 2113 -229
rect 2091 -233 2093 -231
rect 2095 -233 2100 -231
rect 2102 -233 2113 -231
rect 2091 -235 2113 -233
rect 2117 -231 2123 -229
rect 2117 -233 2119 -231
rect 2121 -233 2123 -231
rect 2117 -235 2123 -233
rect 2131 -232 2133 -219
rect 2141 -222 2143 -219
rect 2137 -224 2143 -222
rect 2137 -226 2139 -224
rect 2141 -226 2143 -224
rect 2162 -220 2164 -215
rect 2172 -220 2174 -215
rect 2182 -217 2184 -212
rect 2206 -214 2208 -204
rect 2216 -212 2218 -208
rect 2223 -212 2225 -204
rect 2274 -204 2293 -202
rect 2233 -212 2235 -207
rect 2240 -212 2242 -207
rect 2250 -212 2252 -207
rect 2137 -228 2143 -226
rect 2131 -234 2137 -232
rect 1989 -238 1998 -236
rect 2006 -238 2008 -235
rect 2013 -238 2015 -235
rect 2031 -238 2033 -235
rect 2041 -238 2043 -235
rect 2051 -238 2053 -235
rect 2073 -238 2075 -235
rect 2083 -238 2085 -235
rect 2093 -238 2095 -235
rect 2111 -238 2113 -235
rect 2118 -238 2120 -235
rect 2131 -236 2133 -234
rect 2135 -236 2137 -234
rect 2128 -238 2137 -236
rect 1996 -241 1998 -238
rect 1996 -259 1998 -254
rect 1963 -270 1965 -266
rect 1983 -270 1985 -266
rect 2006 -268 2008 -263
rect 2013 -268 2015 -263
rect 2128 -241 2130 -238
rect 2141 -241 2143 -228
rect 2162 -236 2164 -226
rect 2172 -229 2174 -226
rect 2182 -229 2184 -226
rect 2168 -231 2174 -229
rect 2168 -233 2170 -231
rect 2172 -233 2174 -231
rect 2168 -235 2174 -233
rect 2178 -231 2184 -229
rect 2178 -233 2180 -231
rect 2182 -233 2184 -231
rect 2178 -235 2184 -233
rect 2158 -238 2164 -236
rect 2158 -240 2160 -238
rect 2162 -240 2164 -238
rect 2128 -259 2130 -254
rect 2031 -270 2033 -266
rect 2041 -270 2043 -266
rect 2051 -270 2053 -266
rect 2073 -270 2075 -266
rect 2083 -270 2085 -266
rect 2093 -270 2095 -266
rect 2111 -268 2113 -263
rect 2118 -268 2120 -263
rect 2158 -242 2164 -240
rect 2162 -245 2164 -242
rect 2169 -245 2171 -235
rect 2182 -238 2184 -235
rect 2206 -238 2208 -220
rect 2216 -229 2218 -220
rect 2212 -231 2218 -229
rect 2212 -233 2214 -231
rect 2216 -233 2218 -231
rect 2212 -235 2218 -233
rect 2223 -233 2225 -220
rect 2233 -223 2235 -220
rect 2229 -225 2235 -223
rect 2229 -227 2231 -225
rect 2233 -227 2235 -225
rect 2229 -229 2235 -227
rect 2223 -235 2235 -233
rect 2240 -234 2242 -220
rect 2274 -214 2276 -204
rect 2284 -212 2286 -208
rect 2291 -212 2293 -204
rect 2301 -212 2303 -207
rect 2308 -212 2310 -207
rect 2318 -212 2320 -207
rect 2250 -224 2252 -221
rect 2247 -226 2253 -224
rect 2247 -228 2249 -226
rect 2251 -228 2253 -226
rect 2247 -230 2253 -228
rect 2206 -249 2208 -246
rect 2199 -251 2208 -249
rect 2216 -250 2218 -235
rect 2222 -241 2228 -239
rect 2222 -243 2224 -241
rect 2226 -243 2228 -241
rect 2222 -245 2228 -243
rect 2223 -250 2225 -245
rect 2233 -250 2235 -235
rect 2239 -236 2245 -234
rect 2239 -238 2241 -236
rect 2243 -238 2245 -236
rect 2239 -240 2245 -238
rect 2240 -250 2242 -240
rect 2250 -248 2252 -230
rect 2274 -238 2276 -220
rect 2284 -229 2286 -220
rect 2280 -231 2286 -229
rect 2280 -233 2282 -231
rect 2284 -233 2286 -231
rect 2280 -235 2286 -233
rect 2291 -233 2293 -220
rect 2301 -223 2303 -220
rect 2297 -225 2303 -223
rect 2297 -227 2299 -225
rect 2301 -227 2303 -225
rect 2297 -229 2303 -227
rect 2291 -235 2303 -233
rect 2308 -234 2310 -220
rect 2318 -224 2320 -221
rect 2315 -226 2321 -224
rect 2315 -228 2317 -226
rect 2319 -228 2321 -226
rect 2315 -230 2321 -228
rect 2199 -253 2201 -251
rect 2203 -253 2205 -251
rect 2199 -255 2205 -253
rect 2182 -261 2184 -256
rect 2141 -270 2143 -266
rect 2162 -270 2164 -266
rect 2169 -270 2171 -266
rect 2274 -249 2276 -246
rect 2267 -251 2276 -249
rect 2284 -250 2286 -235
rect 2290 -241 2296 -239
rect 2290 -243 2292 -241
rect 2294 -243 2296 -241
rect 2290 -245 2296 -243
rect 2291 -250 2293 -245
rect 2301 -250 2303 -235
rect 2307 -236 2313 -234
rect 2307 -238 2309 -236
rect 2311 -238 2313 -236
rect 2307 -240 2313 -238
rect 2308 -250 2310 -240
rect 2318 -248 2320 -230
rect 2267 -253 2269 -251
rect 2271 -253 2273 -251
rect 2267 -255 2273 -253
rect 2216 -270 2218 -266
rect 2223 -270 2225 -266
rect 2233 -270 2235 -266
rect 2240 -270 2242 -266
rect 2250 -270 2252 -266
rect 2284 -270 2286 -266
rect 2291 -270 2293 -266
rect 2301 -270 2303 -266
rect 2308 -270 2310 -266
rect 2318 -270 2320 -266
<< ndif >>
rect 10 251 15 256
rect 8 249 15 251
rect 8 247 10 249
rect 12 247 15 249
rect 8 245 15 247
rect 17 245 22 256
rect 24 247 35 256
rect 37 253 42 256
rect 37 251 44 253
rect 50 251 55 256
rect 37 249 40 251
rect 42 249 44 251
rect 37 247 44 249
rect 48 249 55 251
rect 48 247 50 249
rect 52 247 55 249
rect 24 245 33 247
rect 26 239 33 245
rect 48 245 55 247
rect 57 245 62 256
rect 64 247 75 256
rect 77 253 82 256
rect 77 251 84 253
rect 110 251 115 258
rect 77 249 80 251
rect 82 249 84 251
rect 77 247 84 249
rect 88 249 95 251
rect 88 247 90 249
rect 92 247 95 249
rect 64 245 73 247
rect 26 237 29 239
rect 31 237 33 239
rect 26 235 33 237
rect 66 239 73 245
rect 88 245 95 247
rect 66 237 69 239
rect 71 237 73 239
rect 66 235 73 237
rect 90 238 95 245
rect 97 245 105 251
rect 97 243 100 245
rect 102 243 105 245
rect 97 241 105 243
rect 107 248 115 251
rect 107 246 110 248
rect 112 246 115 248
rect 107 244 115 246
rect 117 256 125 258
rect 117 254 120 256
rect 122 254 125 256
rect 117 244 125 254
rect 127 256 134 258
rect 127 254 130 256
rect 132 254 134 256
rect 127 249 134 254
rect 140 251 145 258
rect 127 247 130 249
rect 132 247 134 249
rect 127 244 134 247
rect 138 249 145 251
rect 138 247 140 249
rect 142 247 145 249
rect 138 245 145 247
rect 107 241 112 244
rect 97 238 102 241
rect 140 238 145 245
rect 147 238 152 258
rect 154 252 161 258
rect 189 252 196 258
rect 154 242 163 252
rect 154 240 157 242
rect 159 240 163 242
rect 154 238 163 240
rect 165 249 172 252
rect 165 247 168 249
rect 170 247 172 249
rect 165 245 172 247
rect 178 249 185 252
rect 178 247 180 249
rect 182 247 185 249
rect 178 245 185 247
rect 165 238 170 245
rect 180 238 185 245
rect 187 242 196 252
rect 187 240 191 242
rect 193 240 196 242
rect 187 238 196 240
rect 198 238 203 258
rect 205 251 210 258
rect 216 256 223 258
rect 216 254 218 256
rect 220 254 223 256
rect 205 249 212 251
rect 205 247 208 249
rect 210 247 212 249
rect 205 245 212 247
rect 216 249 223 254
rect 216 247 218 249
rect 220 247 223 249
rect 205 238 210 245
rect 216 244 223 247
rect 225 256 233 258
rect 225 254 228 256
rect 230 254 233 256
rect 225 244 233 254
rect 235 251 240 258
rect 267 252 274 258
rect 276 256 284 258
rect 276 254 279 256
rect 281 254 284 256
rect 276 252 284 254
rect 286 252 294 258
rect 235 248 243 251
rect 235 246 238 248
rect 240 246 243 248
rect 235 244 243 246
rect 238 241 243 244
rect 245 245 253 251
rect 245 243 248 245
rect 250 243 253 245
rect 245 241 253 243
rect 248 238 253 241
rect 255 249 262 251
rect 255 247 258 249
rect 260 247 262 249
rect 255 245 262 247
rect 267 245 272 252
rect 288 249 294 252
rect 296 256 303 258
rect 296 254 299 256
rect 301 254 303 256
rect 296 252 303 254
rect 296 249 301 252
rect 317 251 322 256
rect 315 249 322 251
rect 288 245 292 249
rect 255 238 260 245
rect 267 243 273 245
rect 267 241 269 243
rect 271 241 273 243
rect 267 239 273 241
rect 286 243 292 245
rect 315 247 317 249
rect 319 247 322 249
rect 315 245 322 247
rect 324 245 329 256
rect 331 247 342 256
rect 344 253 349 256
rect 344 251 351 253
rect 377 251 382 258
rect 344 249 347 251
rect 349 249 351 251
rect 344 247 351 249
rect 355 249 362 251
rect 355 247 357 249
rect 359 247 362 249
rect 331 245 340 247
rect 286 241 288 243
rect 290 241 292 243
rect 286 239 292 241
rect 333 239 340 245
rect 355 245 362 247
rect 333 237 336 239
rect 338 237 340 239
rect 333 235 340 237
rect 357 238 362 245
rect 364 245 372 251
rect 364 243 367 245
rect 369 243 372 245
rect 364 241 372 243
rect 374 248 382 251
rect 374 246 377 248
rect 379 246 382 248
rect 374 244 382 246
rect 384 256 392 258
rect 384 254 387 256
rect 389 254 392 256
rect 384 244 392 254
rect 394 256 401 258
rect 394 254 397 256
rect 399 254 401 256
rect 394 249 401 254
rect 407 251 412 258
rect 394 247 397 249
rect 399 247 401 249
rect 394 244 401 247
rect 405 249 412 251
rect 405 247 407 249
rect 409 247 412 249
rect 405 245 412 247
rect 374 241 379 244
rect 364 238 369 241
rect 407 238 412 245
rect 414 238 419 258
rect 421 252 428 258
rect 456 252 463 258
rect 421 242 430 252
rect 421 240 424 242
rect 426 240 430 242
rect 421 238 430 240
rect 432 249 439 252
rect 432 247 435 249
rect 437 247 439 249
rect 432 245 439 247
rect 445 249 452 252
rect 445 247 447 249
rect 449 247 452 249
rect 445 245 452 247
rect 432 238 437 245
rect 447 238 452 245
rect 454 242 463 252
rect 454 240 458 242
rect 460 240 463 242
rect 454 238 463 240
rect 465 238 470 258
rect 472 251 477 258
rect 483 256 490 258
rect 483 254 485 256
rect 487 254 490 256
rect 472 249 479 251
rect 472 247 475 249
rect 477 247 479 249
rect 472 245 479 247
rect 483 249 490 254
rect 483 247 485 249
rect 487 247 490 249
rect 472 238 477 245
rect 483 244 490 247
rect 492 256 500 258
rect 492 254 495 256
rect 497 254 500 256
rect 492 244 500 254
rect 502 251 507 258
rect 534 252 541 258
rect 543 256 551 258
rect 543 254 546 256
rect 548 254 551 256
rect 543 252 551 254
rect 553 252 561 258
rect 502 248 510 251
rect 502 246 505 248
rect 507 246 510 248
rect 502 244 510 246
rect 505 241 510 244
rect 512 245 520 251
rect 512 243 515 245
rect 517 243 520 245
rect 512 241 520 243
rect 515 238 520 241
rect 522 249 529 251
rect 522 247 525 249
rect 527 247 529 249
rect 522 245 529 247
rect 534 245 539 252
rect 555 249 561 252
rect 563 256 570 258
rect 563 254 566 256
rect 568 254 570 256
rect 563 252 570 254
rect 563 249 568 252
rect 584 251 589 256
rect 582 249 589 251
rect 555 245 559 249
rect 522 238 527 245
rect 534 243 540 245
rect 534 241 536 243
rect 538 241 540 243
rect 534 239 540 241
rect 553 243 559 245
rect 582 247 584 249
rect 586 247 589 249
rect 582 245 589 247
rect 591 245 596 256
rect 598 247 609 256
rect 611 253 616 256
rect 611 251 618 253
rect 644 251 649 258
rect 611 249 614 251
rect 616 249 618 251
rect 611 247 618 249
rect 622 249 629 251
rect 622 247 624 249
rect 626 247 629 249
rect 598 245 607 247
rect 553 241 555 243
rect 557 241 559 243
rect 553 239 559 241
rect 600 239 607 245
rect 622 245 629 247
rect 600 237 603 239
rect 605 237 607 239
rect 600 235 607 237
rect 624 238 629 245
rect 631 245 639 251
rect 631 243 634 245
rect 636 243 639 245
rect 631 241 639 243
rect 641 248 649 251
rect 641 246 644 248
rect 646 246 649 248
rect 641 244 649 246
rect 651 256 659 258
rect 651 254 654 256
rect 656 254 659 256
rect 651 244 659 254
rect 661 256 668 258
rect 661 254 664 256
rect 666 254 668 256
rect 661 249 668 254
rect 674 251 679 258
rect 661 247 664 249
rect 666 247 668 249
rect 661 244 668 247
rect 672 249 679 251
rect 672 247 674 249
rect 676 247 679 249
rect 672 245 679 247
rect 641 241 646 244
rect 631 238 636 241
rect 674 238 679 245
rect 681 238 686 258
rect 688 252 695 258
rect 723 252 730 258
rect 688 242 697 252
rect 688 240 691 242
rect 693 240 697 242
rect 688 238 697 240
rect 699 249 706 252
rect 699 247 702 249
rect 704 247 706 249
rect 699 245 706 247
rect 712 249 719 252
rect 712 247 714 249
rect 716 247 719 249
rect 712 245 719 247
rect 699 238 704 245
rect 714 238 719 245
rect 721 242 730 252
rect 721 240 725 242
rect 727 240 730 242
rect 721 238 730 240
rect 732 238 737 258
rect 739 251 744 258
rect 750 256 757 258
rect 750 254 752 256
rect 754 254 757 256
rect 739 249 746 251
rect 739 247 742 249
rect 744 247 746 249
rect 739 245 746 247
rect 750 249 757 254
rect 750 247 752 249
rect 754 247 757 249
rect 739 238 744 245
rect 750 244 757 247
rect 759 256 767 258
rect 759 254 762 256
rect 764 254 767 256
rect 759 244 767 254
rect 769 251 774 258
rect 801 252 808 258
rect 810 256 818 258
rect 810 254 813 256
rect 815 254 818 256
rect 810 252 818 254
rect 820 252 828 258
rect 769 248 777 251
rect 769 246 772 248
rect 774 246 777 248
rect 769 244 777 246
rect 772 241 777 244
rect 779 245 787 251
rect 779 243 782 245
rect 784 243 787 245
rect 779 241 787 243
rect 782 238 787 241
rect 789 249 796 251
rect 789 247 792 249
rect 794 247 796 249
rect 789 245 796 247
rect 801 245 806 252
rect 822 249 828 252
rect 830 256 837 258
rect 830 254 833 256
rect 835 254 837 256
rect 830 252 837 254
rect 830 249 835 252
rect 851 251 856 256
rect 849 249 856 251
rect 822 245 826 249
rect 789 238 794 245
rect 801 243 807 245
rect 801 241 803 243
rect 805 241 807 243
rect 801 239 807 241
rect 820 243 826 245
rect 849 247 851 249
rect 853 247 856 249
rect 849 245 856 247
rect 858 245 863 256
rect 865 247 876 256
rect 878 253 883 256
rect 878 251 885 253
rect 911 251 916 258
rect 878 249 881 251
rect 883 249 885 251
rect 878 247 885 249
rect 889 249 896 251
rect 889 247 891 249
rect 893 247 896 249
rect 865 245 874 247
rect 820 241 822 243
rect 824 241 826 243
rect 820 239 826 241
rect 867 239 874 245
rect 889 245 896 247
rect 867 237 870 239
rect 872 237 874 239
rect 867 235 874 237
rect 891 238 896 245
rect 898 245 906 251
rect 898 243 901 245
rect 903 243 906 245
rect 898 241 906 243
rect 908 248 916 251
rect 908 246 911 248
rect 913 246 916 248
rect 908 244 916 246
rect 918 256 926 258
rect 918 254 921 256
rect 923 254 926 256
rect 918 244 926 254
rect 928 256 935 258
rect 928 254 931 256
rect 933 254 935 256
rect 928 249 935 254
rect 941 251 946 258
rect 928 247 931 249
rect 933 247 935 249
rect 928 244 935 247
rect 939 249 946 251
rect 939 247 941 249
rect 943 247 946 249
rect 939 245 946 247
rect 908 241 913 244
rect 898 238 903 241
rect 941 238 946 245
rect 948 238 953 258
rect 955 252 962 258
rect 990 252 997 258
rect 955 242 964 252
rect 955 240 958 242
rect 960 240 964 242
rect 955 238 964 240
rect 966 249 973 252
rect 966 247 969 249
rect 971 247 973 249
rect 966 245 973 247
rect 979 249 986 252
rect 979 247 981 249
rect 983 247 986 249
rect 979 245 986 247
rect 966 238 971 245
rect 981 238 986 245
rect 988 242 997 252
rect 988 240 992 242
rect 994 240 997 242
rect 988 238 997 240
rect 999 238 1004 258
rect 1006 251 1011 258
rect 1017 256 1024 258
rect 1017 254 1019 256
rect 1021 254 1024 256
rect 1006 249 1013 251
rect 1006 247 1009 249
rect 1011 247 1013 249
rect 1006 245 1013 247
rect 1017 249 1024 254
rect 1017 247 1019 249
rect 1021 247 1024 249
rect 1006 238 1011 245
rect 1017 244 1024 247
rect 1026 256 1034 258
rect 1026 254 1029 256
rect 1031 254 1034 256
rect 1026 244 1034 254
rect 1036 251 1041 258
rect 1068 252 1075 258
rect 1077 256 1085 258
rect 1077 254 1080 256
rect 1082 254 1085 256
rect 1077 252 1085 254
rect 1087 252 1095 258
rect 1036 248 1044 251
rect 1036 246 1039 248
rect 1041 246 1044 248
rect 1036 244 1044 246
rect 1039 241 1044 244
rect 1046 245 1054 251
rect 1046 243 1049 245
rect 1051 243 1054 245
rect 1046 241 1054 243
rect 1049 238 1054 241
rect 1056 249 1063 251
rect 1056 247 1059 249
rect 1061 247 1063 249
rect 1056 245 1063 247
rect 1068 245 1073 252
rect 1089 249 1095 252
rect 1097 256 1104 258
rect 1097 254 1100 256
rect 1102 254 1104 256
rect 1097 252 1104 254
rect 1097 249 1102 252
rect 1118 251 1123 256
rect 1116 249 1123 251
rect 1089 245 1093 249
rect 1056 238 1061 245
rect 1068 243 1074 245
rect 1068 241 1070 243
rect 1072 241 1074 243
rect 1068 239 1074 241
rect 1087 243 1093 245
rect 1116 247 1118 249
rect 1120 247 1123 249
rect 1116 245 1123 247
rect 1125 245 1130 256
rect 1132 247 1143 256
rect 1145 253 1150 256
rect 1145 251 1152 253
rect 1178 251 1183 258
rect 1145 249 1148 251
rect 1150 249 1152 251
rect 1145 247 1152 249
rect 1156 249 1163 251
rect 1156 247 1158 249
rect 1160 247 1163 249
rect 1132 245 1141 247
rect 1087 241 1089 243
rect 1091 241 1093 243
rect 1087 239 1093 241
rect 1134 239 1141 245
rect 1156 245 1163 247
rect 1134 237 1137 239
rect 1139 237 1141 239
rect 1134 235 1141 237
rect 1158 238 1163 245
rect 1165 245 1173 251
rect 1165 243 1168 245
rect 1170 243 1173 245
rect 1165 241 1173 243
rect 1175 248 1183 251
rect 1175 246 1178 248
rect 1180 246 1183 248
rect 1175 244 1183 246
rect 1185 256 1193 258
rect 1185 254 1188 256
rect 1190 254 1193 256
rect 1185 244 1193 254
rect 1195 256 1202 258
rect 1195 254 1198 256
rect 1200 254 1202 256
rect 1195 249 1202 254
rect 1208 251 1213 258
rect 1195 247 1198 249
rect 1200 247 1202 249
rect 1195 244 1202 247
rect 1206 249 1213 251
rect 1206 247 1208 249
rect 1210 247 1213 249
rect 1206 245 1213 247
rect 1175 241 1180 244
rect 1165 238 1170 241
rect 1208 238 1213 245
rect 1215 238 1220 258
rect 1222 252 1229 258
rect 1257 252 1264 258
rect 1222 242 1231 252
rect 1222 240 1225 242
rect 1227 240 1231 242
rect 1222 238 1231 240
rect 1233 249 1240 252
rect 1233 247 1236 249
rect 1238 247 1240 249
rect 1233 245 1240 247
rect 1246 249 1253 252
rect 1246 247 1248 249
rect 1250 247 1253 249
rect 1246 245 1253 247
rect 1233 238 1238 245
rect 1248 238 1253 245
rect 1255 242 1264 252
rect 1255 240 1259 242
rect 1261 240 1264 242
rect 1255 238 1264 240
rect 1266 238 1271 258
rect 1273 251 1278 258
rect 1284 256 1291 258
rect 1284 254 1286 256
rect 1288 254 1291 256
rect 1273 249 1280 251
rect 1273 247 1276 249
rect 1278 247 1280 249
rect 1273 245 1280 247
rect 1284 249 1291 254
rect 1284 247 1286 249
rect 1288 247 1291 249
rect 1273 238 1278 245
rect 1284 244 1291 247
rect 1293 256 1301 258
rect 1293 254 1296 256
rect 1298 254 1301 256
rect 1293 244 1301 254
rect 1303 251 1308 258
rect 1335 252 1342 258
rect 1344 256 1352 258
rect 1344 254 1347 256
rect 1349 254 1352 256
rect 1344 252 1352 254
rect 1354 252 1362 258
rect 1303 248 1311 251
rect 1303 246 1306 248
rect 1308 246 1311 248
rect 1303 244 1311 246
rect 1306 241 1311 244
rect 1313 245 1321 251
rect 1313 243 1316 245
rect 1318 243 1321 245
rect 1313 241 1321 243
rect 1316 238 1321 241
rect 1323 249 1330 251
rect 1323 247 1326 249
rect 1328 247 1330 249
rect 1323 245 1330 247
rect 1335 245 1340 252
rect 1356 249 1362 252
rect 1364 256 1371 258
rect 1364 254 1367 256
rect 1369 254 1371 256
rect 1364 252 1371 254
rect 1364 249 1369 252
rect 1385 251 1390 256
rect 1383 249 1390 251
rect 1356 245 1360 249
rect 1323 238 1328 245
rect 1335 243 1341 245
rect 1335 241 1337 243
rect 1339 241 1341 243
rect 1335 239 1341 241
rect 1354 243 1360 245
rect 1383 247 1385 249
rect 1387 247 1390 249
rect 1383 245 1390 247
rect 1392 245 1397 256
rect 1399 247 1410 256
rect 1412 253 1417 256
rect 1412 251 1419 253
rect 1445 251 1450 258
rect 1412 249 1415 251
rect 1417 249 1419 251
rect 1412 247 1419 249
rect 1423 249 1430 251
rect 1423 247 1425 249
rect 1427 247 1430 249
rect 1399 245 1408 247
rect 1354 241 1356 243
rect 1358 241 1360 243
rect 1354 239 1360 241
rect 1401 239 1408 245
rect 1423 245 1430 247
rect 1401 237 1404 239
rect 1406 237 1408 239
rect 1401 235 1408 237
rect 1425 238 1430 245
rect 1432 245 1440 251
rect 1432 243 1435 245
rect 1437 243 1440 245
rect 1432 241 1440 243
rect 1442 248 1450 251
rect 1442 246 1445 248
rect 1447 246 1450 248
rect 1442 244 1450 246
rect 1452 256 1460 258
rect 1452 254 1455 256
rect 1457 254 1460 256
rect 1452 244 1460 254
rect 1462 256 1469 258
rect 1462 254 1465 256
rect 1467 254 1469 256
rect 1462 249 1469 254
rect 1475 251 1480 258
rect 1462 247 1465 249
rect 1467 247 1469 249
rect 1462 244 1469 247
rect 1473 249 1480 251
rect 1473 247 1475 249
rect 1477 247 1480 249
rect 1473 245 1480 247
rect 1442 241 1447 244
rect 1432 238 1437 241
rect 1475 238 1480 245
rect 1482 238 1487 258
rect 1489 252 1496 258
rect 1524 252 1531 258
rect 1489 242 1498 252
rect 1489 240 1492 242
rect 1494 240 1498 242
rect 1489 238 1498 240
rect 1500 249 1507 252
rect 1500 247 1503 249
rect 1505 247 1507 249
rect 1500 245 1507 247
rect 1513 249 1520 252
rect 1513 247 1515 249
rect 1517 247 1520 249
rect 1513 245 1520 247
rect 1500 238 1505 245
rect 1515 238 1520 245
rect 1522 242 1531 252
rect 1522 240 1526 242
rect 1528 240 1531 242
rect 1522 238 1531 240
rect 1533 238 1538 258
rect 1540 251 1545 258
rect 1551 256 1558 258
rect 1551 254 1553 256
rect 1555 254 1558 256
rect 1540 249 1547 251
rect 1540 247 1543 249
rect 1545 247 1547 249
rect 1540 245 1547 247
rect 1551 249 1558 254
rect 1551 247 1553 249
rect 1555 247 1558 249
rect 1540 238 1545 245
rect 1551 244 1558 247
rect 1560 256 1568 258
rect 1560 254 1563 256
rect 1565 254 1568 256
rect 1560 244 1568 254
rect 1570 251 1575 258
rect 1602 252 1609 258
rect 1611 256 1619 258
rect 1611 254 1614 256
rect 1616 254 1619 256
rect 1611 252 1619 254
rect 1621 252 1629 258
rect 1570 248 1578 251
rect 1570 246 1573 248
rect 1575 246 1578 248
rect 1570 244 1578 246
rect 1573 241 1578 244
rect 1580 245 1588 251
rect 1580 243 1583 245
rect 1585 243 1588 245
rect 1580 241 1588 243
rect 1583 238 1588 241
rect 1590 249 1597 251
rect 1590 247 1593 249
rect 1595 247 1597 249
rect 1590 245 1597 247
rect 1602 245 1607 252
rect 1623 249 1629 252
rect 1631 256 1638 258
rect 1631 254 1634 256
rect 1636 254 1638 256
rect 1631 252 1638 254
rect 1631 249 1636 252
rect 1652 251 1657 256
rect 1650 249 1657 251
rect 1623 245 1627 249
rect 1590 238 1595 245
rect 1602 243 1608 245
rect 1602 241 1604 243
rect 1606 241 1608 243
rect 1602 239 1608 241
rect 1621 243 1627 245
rect 1650 247 1652 249
rect 1654 247 1657 249
rect 1650 245 1657 247
rect 1659 245 1664 256
rect 1666 247 1677 256
rect 1679 253 1684 256
rect 1679 251 1686 253
rect 1712 251 1717 258
rect 1679 249 1682 251
rect 1684 249 1686 251
rect 1679 247 1686 249
rect 1690 249 1697 251
rect 1690 247 1692 249
rect 1694 247 1697 249
rect 1666 245 1675 247
rect 1621 241 1623 243
rect 1625 241 1627 243
rect 1621 239 1627 241
rect 1668 239 1675 245
rect 1690 245 1697 247
rect 1668 237 1671 239
rect 1673 237 1675 239
rect 1668 235 1675 237
rect 1692 238 1697 245
rect 1699 245 1707 251
rect 1699 243 1702 245
rect 1704 243 1707 245
rect 1699 241 1707 243
rect 1709 248 1717 251
rect 1709 246 1712 248
rect 1714 246 1717 248
rect 1709 244 1717 246
rect 1719 256 1727 258
rect 1719 254 1722 256
rect 1724 254 1727 256
rect 1719 244 1727 254
rect 1729 256 1736 258
rect 1729 254 1732 256
rect 1734 254 1736 256
rect 1729 249 1736 254
rect 1742 251 1747 258
rect 1729 247 1732 249
rect 1734 247 1736 249
rect 1729 244 1736 247
rect 1740 249 1747 251
rect 1740 247 1742 249
rect 1744 247 1747 249
rect 1740 245 1747 247
rect 1709 241 1714 244
rect 1699 238 1704 241
rect 1742 238 1747 245
rect 1749 238 1754 258
rect 1756 252 1763 258
rect 1791 252 1798 258
rect 1756 242 1765 252
rect 1756 240 1759 242
rect 1761 240 1765 242
rect 1756 238 1765 240
rect 1767 249 1774 252
rect 1767 247 1770 249
rect 1772 247 1774 249
rect 1767 245 1774 247
rect 1780 249 1787 252
rect 1780 247 1782 249
rect 1784 247 1787 249
rect 1780 245 1787 247
rect 1767 238 1772 245
rect 1782 238 1787 245
rect 1789 242 1798 252
rect 1789 240 1793 242
rect 1795 240 1798 242
rect 1789 238 1798 240
rect 1800 238 1805 258
rect 1807 251 1812 258
rect 1818 256 1825 258
rect 1818 254 1820 256
rect 1822 254 1825 256
rect 1807 249 1814 251
rect 1807 247 1810 249
rect 1812 247 1814 249
rect 1807 245 1814 247
rect 1818 249 1825 254
rect 1818 247 1820 249
rect 1822 247 1825 249
rect 1807 238 1812 245
rect 1818 244 1825 247
rect 1827 256 1835 258
rect 1827 254 1830 256
rect 1832 254 1835 256
rect 1827 244 1835 254
rect 1837 251 1842 258
rect 1869 252 1876 258
rect 1878 256 1886 258
rect 1878 254 1881 256
rect 1883 254 1886 256
rect 1878 252 1886 254
rect 1888 252 1896 258
rect 1837 248 1845 251
rect 1837 246 1840 248
rect 1842 246 1845 248
rect 1837 244 1845 246
rect 1840 241 1845 244
rect 1847 245 1855 251
rect 1847 243 1850 245
rect 1852 243 1855 245
rect 1847 241 1855 243
rect 1850 238 1855 241
rect 1857 249 1864 251
rect 1857 247 1860 249
rect 1862 247 1864 249
rect 1857 245 1864 247
rect 1869 245 1874 252
rect 1890 249 1896 252
rect 1898 256 1905 258
rect 1898 254 1901 256
rect 1903 254 1905 256
rect 1898 252 1905 254
rect 1912 256 1919 258
rect 1912 254 1914 256
rect 1916 254 1919 256
rect 1912 252 1919 254
rect 1898 249 1903 252
rect 1914 249 1919 252
rect 1921 253 1926 258
rect 1921 249 1935 253
rect 1890 245 1894 249
rect 1857 238 1862 245
rect 1869 243 1875 245
rect 1869 241 1871 243
rect 1873 241 1875 243
rect 1869 239 1875 241
rect 1888 243 1894 245
rect 1926 248 1935 249
rect 1926 246 1928 248
rect 1930 246 1935 248
rect 1926 244 1935 246
rect 1937 251 1945 253
rect 1937 249 1940 251
rect 1942 249 1945 251
rect 1937 244 1945 249
rect 1947 249 1955 253
rect 1947 247 1950 249
rect 1952 247 1955 249
rect 1947 244 1955 247
rect 1888 241 1890 243
rect 1892 241 1894 243
rect 1888 239 1894 241
rect 1950 241 1955 244
rect 1957 241 1962 253
rect 1964 241 1972 253
rect 1998 251 2003 258
rect 1976 249 1983 251
rect 1976 247 1978 249
rect 1980 247 1983 249
rect 1976 245 1983 247
rect 1966 239 1972 241
rect 1966 237 1968 239
rect 1970 237 1972 239
rect 1978 238 1983 245
rect 1985 245 1993 251
rect 1985 243 1988 245
rect 1990 243 1993 245
rect 1985 241 1993 243
rect 1995 248 2003 251
rect 1995 246 1998 248
rect 2000 246 2003 248
rect 1995 244 2003 246
rect 2005 256 2013 258
rect 2005 254 2008 256
rect 2010 254 2013 256
rect 2005 244 2013 254
rect 2015 256 2022 258
rect 2015 254 2018 256
rect 2020 254 2022 256
rect 2015 249 2022 254
rect 2028 251 2033 258
rect 2015 247 2018 249
rect 2020 247 2022 249
rect 2015 244 2022 247
rect 2026 249 2033 251
rect 2026 247 2028 249
rect 2030 247 2033 249
rect 2026 245 2033 247
rect 1995 241 2000 244
rect 1985 238 1990 241
rect 1966 235 1972 237
rect 2028 238 2033 245
rect 2035 238 2040 258
rect 2042 252 2049 258
rect 2077 252 2084 258
rect 2042 242 2051 252
rect 2042 240 2045 242
rect 2047 240 2051 242
rect 2042 238 2051 240
rect 2053 249 2060 252
rect 2053 247 2056 249
rect 2058 247 2060 249
rect 2053 245 2060 247
rect 2066 249 2073 252
rect 2066 247 2068 249
rect 2070 247 2073 249
rect 2066 245 2073 247
rect 2053 238 2058 245
rect 2068 238 2073 245
rect 2075 242 2084 252
rect 2075 240 2079 242
rect 2081 240 2084 242
rect 2075 238 2084 240
rect 2086 238 2091 258
rect 2093 251 2098 258
rect 2104 256 2111 258
rect 2104 254 2106 256
rect 2108 254 2111 256
rect 2093 249 2100 251
rect 2093 247 2096 249
rect 2098 247 2100 249
rect 2093 245 2100 247
rect 2104 249 2111 254
rect 2104 247 2106 249
rect 2108 247 2111 249
rect 2093 238 2098 245
rect 2104 244 2111 247
rect 2113 256 2121 258
rect 2113 254 2116 256
rect 2118 254 2121 256
rect 2113 244 2121 254
rect 2123 251 2128 258
rect 2155 252 2162 258
rect 2164 256 2172 258
rect 2164 254 2167 256
rect 2169 254 2172 256
rect 2164 252 2172 254
rect 2174 252 2182 258
rect 2123 248 2131 251
rect 2123 246 2126 248
rect 2128 246 2131 248
rect 2123 244 2131 246
rect 2126 241 2131 244
rect 2133 245 2141 251
rect 2133 243 2136 245
rect 2138 243 2141 245
rect 2133 241 2141 243
rect 2136 238 2141 241
rect 2143 249 2150 251
rect 2143 247 2146 249
rect 2148 247 2150 249
rect 2143 245 2150 247
rect 2155 245 2160 252
rect 2176 249 2182 252
rect 2184 256 2191 258
rect 2184 254 2187 256
rect 2189 254 2191 256
rect 2184 252 2191 254
rect 2245 252 2250 253
rect 2184 249 2189 252
rect 2199 250 2206 252
rect 2176 245 2180 249
rect 2143 238 2148 245
rect 2155 243 2161 245
rect 2155 241 2157 243
rect 2159 241 2161 243
rect 2155 239 2161 241
rect 2174 243 2180 245
rect 2199 248 2201 250
rect 2203 248 2206 250
rect 2199 246 2206 248
rect 2208 250 2216 252
rect 2208 248 2211 250
rect 2213 248 2216 250
rect 2208 246 2216 248
rect 2174 241 2176 243
rect 2178 241 2180 243
rect 2174 239 2180 241
rect 2210 244 2216 246
rect 2218 244 2223 252
rect 2225 248 2233 252
rect 2225 246 2228 248
rect 2230 246 2233 248
rect 2225 244 2233 246
rect 2235 244 2240 252
rect 2242 248 2250 252
rect 2242 246 2245 248
rect 2247 246 2250 248
rect 2242 244 2250 246
rect 2252 251 2259 253
rect 2313 252 2318 253
rect 2252 249 2255 251
rect 2257 249 2259 251
rect 2252 247 2259 249
rect 2267 250 2274 252
rect 2267 248 2269 250
rect 2271 248 2274 250
rect 2252 244 2257 247
rect 2267 246 2274 248
rect 2276 250 2284 252
rect 2276 248 2279 250
rect 2281 248 2284 250
rect 2276 246 2284 248
rect 2278 244 2284 246
rect 2286 244 2291 252
rect 2293 248 2301 252
rect 2293 246 2296 248
rect 2298 246 2301 248
rect 2293 244 2301 246
rect 2303 244 2308 252
rect 2310 248 2318 252
rect 2310 246 2313 248
rect 2315 246 2318 248
rect 2310 244 2318 246
rect 2320 251 2327 253
rect 2320 249 2323 251
rect 2325 249 2327 251
rect 2320 247 2327 249
rect 2320 244 2325 247
rect 26 227 33 229
rect 26 225 29 227
rect 31 225 33 227
rect 26 219 33 225
rect 66 227 73 229
rect 66 225 69 227
rect 71 225 73 227
rect 8 217 15 219
rect 8 215 10 217
rect 12 215 15 217
rect 8 213 15 215
rect 10 208 15 213
rect 17 208 22 219
rect 24 217 33 219
rect 66 219 73 225
rect 48 217 55 219
rect 24 208 35 217
rect 37 215 44 217
rect 37 213 40 215
rect 42 213 44 215
rect 48 215 50 217
rect 52 215 55 217
rect 48 213 55 215
rect 37 211 44 213
rect 37 208 42 211
rect 50 208 55 213
rect 57 208 62 219
rect 64 217 73 219
rect 90 219 95 226
rect 88 217 95 219
rect 64 208 75 217
rect 77 215 84 217
rect 77 213 80 215
rect 82 213 84 215
rect 88 215 90 217
rect 92 215 95 217
rect 88 213 95 215
rect 97 223 102 226
rect 97 221 105 223
rect 97 219 100 221
rect 102 219 105 221
rect 97 213 105 219
rect 107 220 112 223
rect 107 218 115 220
rect 107 216 110 218
rect 112 216 115 218
rect 107 213 115 216
rect 77 211 84 213
rect 77 208 82 211
rect 110 206 115 213
rect 117 210 125 220
rect 117 208 120 210
rect 122 208 125 210
rect 117 206 125 208
rect 127 217 134 220
rect 140 219 145 226
rect 127 215 130 217
rect 132 215 134 217
rect 127 210 134 215
rect 138 217 145 219
rect 138 215 140 217
rect 142 215 145 217
rect 138 213 145 215
rect 127 208 130 210
rect 132 208 134 210
rect 127 206 134 208
rect 140 206 145 213
rect 147 206 152 226
rect 154 224 163 226
rect 154 222 157 224
rect 159 222 163 224
rect 154 212 163 222
rect 165 219 170 226
rect 180 219 185 226
rect 165 217 172 219
rect 165 215 168 217
rect 170 215 172 217
rect 165 212 172 215
rect 178 217 185 219
rect 178 215 180 217
rect 182 215 185 217
rect 178 212 185 215
rect 187 224 196 226
rect 187 222 191 224
rect 193 222 196 224
rect 187 212 196 222
rect 154 206 161 212
rect 189 206 196 212
rect 198 206 203 226
rect 205 219 210 226
rect 248 223 253 226
rect 238 220 243 223
rect 205 217 212 219
rect 205 215 208 217
rect 210 215 212 217
rect 205 213 212 215
rect 216 217 223 220
rect 216 215 218 217
rect 220 215 223 217
rect 205 206 210 213
rect 216 210 223 215
rect 216 208 218 210
rect 220 208 223 210
rect 216 206 223 208
rect 225 210 233 220
rect 225 208 228 210
rect 230 208 233 210
rect 225 206 233 208
rect 235 218 243 220
rect 235 216 238 218
rect 240 216 243 218
rect 235 213 243 216
rect 245 221 253 223
rect 245 219 248 221
rect 250 219 253 221
rect 245 213 253 219
rect 255 219 260 226
rect 267 223 273 225
rect 267 221 269 223
rect 271 221 273 223
rect 267 219 273 221
rect 286 223 292 225
rect 333 227 340 229
rect 333 225 336 227
rect 338 225 340 227
rect 286 221 288 223
rect 290 221 292 223
rect 286 219 292 221
rect 255 217 262 219
rect 255 215 258 217
rect 260 215 262 217
rect 255 213 262 215
rect 235 206 240 213
rect 267 212 272 219
rect 288 215 292 219
rect 333 219 340 225
rect 315 217 322 219
rect 315 215 317 217
rect 319 215 322 217
rect 288 212 294 215
rect 267 206 274 212
rect 276 210 284 212
rect 276 208 279 210
rect 281 208 284 210
rect 276 206 284 208
rect 286 206 294 212
rect 296 212 301 215
rect 315 213 322 215
rect 296 210 303 212
rect 296 208 299 210
rect 301 208 303 210
rect 317 208 322 213
rect 324 208 329 219
rect 331 217 340 219
rect 357 219 362 226
rect 355 217 362 219
rect 331 208 342 217
rect 344 215 351 217
rect 344 213 347 215
rect 349 213 351 215
rect 355 215 357 217
rect 359 215 362 217
rect 355 213 362 215
rect 364 223 369 226
rect 364 221 372 223
rect 364 219 367 221
rect 369 219 372 221
rect 364 213 372 219
rect 374 220 379 223
rect 374 218 382 220
rect 374 216 377 218
rect 379 216 382 218
rect 374 213 382 216
rect 344 211 351 213
rect 344 208 349 211
rect 296 206 303 208
rect 377 206 382 213
rect 384 210 392 220
rect 384 208 387 210
rect 389 208 392 210
rect 384 206 392 208
rect 394 217 401 220
rect 407 219 412 226
rect 394 215 397 217
rect 399 215 401 217
rect 394 210 401 215
rect 405 217 412 219
rect 405 215 407 217
rect 409 215 412 217
rect 405 213 412 215
rect 394 208 397 210
rect 399 208 401 210
rect 394 206 401 208
rect 407 206 412 213
rect 414 206 419 226
rect 421 224 430 226
rect 421 222 424 224
rect 426 222 430 224
rect 421 212 430 222
rect 432 219 437 226
rect 447 219 452 226
rect 432 217 439 219
rect 432 215 435 217
rect 437 215 439 217
rect 432 212 439 215
rect 445 217 452 219
rect 445 215 447 217
rect 449 215 452 217
rect 445 212 452 215
rect 454 224 463 226
rect 454 222 458 224
rect 460 222 463 224
rect 454 212 463 222
rect 421 206 428 212
rect 456 206 463 212
rect 465 206 470 226
rect 472 219 477 226
rect 515 223 520 226
rect 505 220 510 223
rect 472 217 479 219
rect 472 215 475 217
rect 477 215 479 217
rect 472 213 479 215
rect 483 217 490 220
rect 483 215 485 217
rect 487 215 490 217
rect 472 206 477 213
rect 483 210 490 215
rect 483 208 485 210
rect 487 208 490 210
rect 483 206 490 208
rect 492 210 500 220
rect 492 208 495 210
rect 497 208 500 210
rect 492 206 500 208
rect 502 218 510 220
rect 502 216 505 218
rect 507 216 510 218
rect 502 213 510 216
rect 512 221 520 223
rect 512 219 515 221
rect 517 219 520 221
rect 512 213 520 219
rect 522 219 527 226
rect 534 223 540 225
rect 534 221 536 223
rect 538 221 540 223
rect 534 219 540 221
rect 553 223 559 225
rect 600 227 607 229
rect 600 225 603 227
rect 605 225 607 227
rect 553 221 555 223
rect 557 221 559 223
rect 553 219 559 221
rect 522 217 529 219
rect 522 215 525 217
rect 527 215 529 217
rect 522 213 529 215
rect 502 206 507 213
rect 534 212 539 219
rect 555 215 559 219
rect 600 219 607 225
rect 582 217 589 219
rect 582 215 584 217
rect 586 215 589 217
rect 555 212 561 215
rect 534 206 541 212
rect 543 210 551 212
rect 543 208 546 210
rect 548 208 551 210
rect 543 206 551 208
rect 553 206 561 212
rect 563 212 568 215
rect 582 213 589 215
rect 563 210 570 212
rect 563 208 566 210
rect 568 208 570 210
rect 584 208 589 213
rect 591 208 596 219
rect 598 217 607 219
rect 624 219 629 226
rect 622 217 629 219
rect 598 208 609 217
rect 611 215 618 217
rect 611 213 614 215
rect 616 213 618 215
rect 622 215 624 217
rect 626 215 629 217
rect 622 213 629 215
rect 631 223 636 226
rect 631 221 639 223
rect 631 219 634 221
rect 636 219 639 221
rect 631 213 639 219
rect 641 220 646 223
rect 641 218 649 220
rect 641 216 644 218
rect 646 216 649 218
rect 641 213 649 216
rect 611 211 618 213
rect 611 208 616 211
rect 563 206 570 208
rect 644 206 649 213
rect 651 210 659 220
rect 651 208 654 210
rect 656 208 659 210
rect 651 206 659 208
rect 661 217 668 220
rect 674 219 679 226
rect 661 215 664 217
rect 666 215 668 217
rect 661 210 668 215
rect 672 217 679 219
rect 672 215 674 217
rect 676 215 679 217
rect 672 213 679 215
rect 661 208 664 210
rect 666 208 668 210
rect 661 206 668 208
rect 674 206 679 213
rect 681 206 686 226
rect 688 224 697 226
rect 688 222 691 224
rect 693 222 697 224
rect 688 212 697 222
rect 699 219 704 226
rect 714 219 719 226
rect 699 217 706 219
rect 699 215 702 217
rect 704 215 706 217
rect 699 212 706 215
rect 712 217 719 219
rect 712 215 714 217
rect 716 215 719 217
rect 712 212 719 215
rect 721 224 730 226
rect 721 222 725 224
rect 727 222 730 224
rect 721 212 730 222
rect 688 206 695 212
rect 723 206 730 212
rect 732 206 737 226
rect 739 219 744 226
rect 782 223 787 226
rect 772 220 777 223
rect 739 217 746 219
rect 739 215 742 217
rect 744 215 746 217
rect 739 213 746 215
rect 750 217 757 220
rect 750 215 752 217
rect 754 215 757 217
rect 739 206 744 213
rect 750 210 757 215
rect 750 208 752 210
rect 754 208 757 210
rect 750 206 757 208
rect 759 210 767 220
rect 759 208 762 210
rect 764 208 767 210
rect 759 206 767 208
rect 769 218 777 220
rect 769 216 772 218
rect 774 216 777 218
rect 769 213 777 216
rect 779 221 787 223
rect 779 219 782 221
rect 784 219 787 221
rect 779 213 787 219
rect 789 219 794 226
rect 801 223 807 225
rect 801 221 803 223
rect 805 221 807 223
rect 801 219 807 221
rect 820 223 826 225
rect 867 227 874 229
rect 867 225 870 227
rect 872 225 874 227
rect 820 221 822 223
rect 824 221 826 223
rect 820 219 826 221
rect 789 217 796 219
rect 789 215 792 217
rect 794 215 796 217
rect 789 213 796 215
rect 769 206 774 213
rect 801 212 806 219
rect 822 215 826 219
rect 867 219 874 225
rect 849 217 856 219
rect 849 215 851 217
rect 853 215 856 217
rect 822 212 828 215
rect 801 206 808 212
rect 810 210 818 212
rect 810 208 813 210
rect 815 208 818 210
rect 810 206 818 208
rect 820 206 828 212
rect 830 212 835 215
rect 849 213 856 215
rect 830 210 837 212
rect 830 208 833 210
rect 835 208 837 210
rect 851 208 856 213
rect 858 208 863 219
rect 865 217 874 219
rect 891 219 896 226
rect 889 217 896 219
rect 865 208 876 217
rect 878 215 885 217
rect 878 213 881 215
rect 883 213 885 215
rect 889 215 891 217
rect 893 215 896 217
rect 889 213 896 215
rect 898 223 903 226
rect 898 221 906 223
rect 898 219 901 221
rect 903 219 906 221
rect 898 213 906 219
rect 908 220 913 223
rect 908 218 916 220
rect 908 216 911 218
rect 913 216 916 218
rect 908 213 916 216
rect 878 211 885 213
rect 878 208 883 211
rect 830 206 837 208
rect 911 206 916 213
rect 918 210 926 220
rect 918 208 921 210
rect 923 208 926 210
rect 918 206 926 208
rect 928 217 935 220
rect 941 219 946 226
rect 928 215 931 217
rect 933 215 935 217
rect 928 210 935 215
rect 939 217 946 219
rect 939 215 941 217
rect 943 215 946 217
rect 939 213 946 215
rect 928 208 931 210
rect 933 208 935 210
rect 928 206 935 208
rect 941 206 946 213
rect 948 206 953 226
rect 955 224 964 226
rect 955 222 958 224
rect 960 222 964 224
rect 955 212 964 222
rect 966 219 971 226
rect 981 219 986 226
rect 966 217 973 219
rect 966 215 969 217
rect 971 215 973 217
rect 966 212 973 215
rect 979 217 986 219
rect 979 215 981 217
rect 983 215 986 217
rect 979 212 986 215
rect 988 224 997 226
rect 988 222 992 224
rect 994 222 997 224
rect 988 212 997 222
rect 955 206 962 212
rect 990 206 997 212
rect 999 206 1004 226
rect 1006 219 1011 226
rect 1049 223 1054 226
rect 1039 220 1044 223
rect 1006 217 1013 219
rect 1006 215 1009 217
rect 1011 215 1013 217
rect 1006 213 1013 215
rect 1017 217 1024 220
rect 1017 215 1019 217
rect 1021 215 1024 217
rect 1006 206 1011 213
rect 1017 210 1024 215
rect 1017 208 1019 210
rect 1021 208 1024 210
rect 1017 206 1024 208
rect 1026 210 1034 220
rect 1026 208 1029 210
rect 1031 208 1034 210
rect 1026 206 1034 208
rect 1036 218 1044 220
rect 1036 216 1039 218
rect 1041 216 1044 218
rect 1036 213 1044 216
rect 1046 221 1054 223
rect 1046 219 1049 221
rect 1051 219 1054 221
rect 1046 213 1054 219
rect 1056 219 1061 226
rect 1068 223 1074 225
rect 1068 221 1070 223
rect 1072 221 1074 223
rect 1068 219 1074 221
rect 1087 223 1093 225
rect 1134 227 1141 229
rect 1134 225 1137 227
rect 1139 225 1141 227
rect 1087 221 1089 223
rect 1091 221 1093 223
rect 1087 219 1093 221
rect 1056 217 1063 219
rect 1056 215 1059 217
rect 1061 215 1063 217
rect 1056 213 1063 215
rect 1036 206 1041 213
rect 1068 212 1073 219
rect 1089 215 1093 219
rect 1134 219 1141 225
rect 1116 217 1123 219
rect 1116 215 1118 217
rect 1120 215 1123 217
rect 1089 212 1095 215
rect 1068 206 1075 212
rect 1077 210 1085 212
rect 1077 208 1080 210
rect 1082 208 1085 210
rect 1077 206 1085 208
rect 1087 206 1095 212
rect 1097 212 1102 215
rect 1116 213 1123 215
rect 1097 210 1104 212
rect 1097 208 1100 210
rect 1102 208 1104 210
rect 1118 208 1123 213
rect 1125 208 1130 219
rect 1132 217 1141 219
rect 1158 219 1163 226
rect 1156 217 1163 219
rect 1132 208 1143 217
rect 1145 215 1152 217
rect 1145 213 1148 215
rect 1150 213 1152 215
rect 1156 215 1158 217
rect 1160 215 1163 217
rect 1156 213 1163 215
rect 1165 223 1170 226
rect 1165 221 1173 223
rect 1165 219 1168 221
rect 1170 219 1173 221
rect 1165 213 1173 219
rect 1175 220 1180 223
rect 1175 218 1183 220
rect 1175 216 1178 218
rect 1180 216 1183 218
rect 1175 213 1183 216
rect 1145 211 1152 213
rect 1145 208 1150 211
rect 1097 206 1104 208
rect 1178 206 1183 213
rect 1185 210 1193 220
rect 1185 208 1188 210
rect 1190 208 1193 210
rect 1185 206 1193 208
rect 1195 217 1202 220
rect 1208 219 1213 226
rect 1195 215 1198 217
rect 1200 215 1202 217
rect 1195 210 1202 215
rect 1206 217 1213 219
rect 1206 215 1208 217
rect 1210 215 1213 217
rect 1206 213 1213 215
rect 1195 208 1198 210
rect 1200 208 1202 210
rect 1195 206 1202 208
rect 1208 206 1213 213
rect 1215 206 1220 226
rect 1222 224 1231 226
rect 1222 222 1225 224
rect 1227 222 1231 224
rect 1222 212 1231 222
rect 1233 219 1238 226
rect 1248 219 1253 226
rect 1233 217 1240 219
rect 1233 215 1236 217
rect 1238 215 1240 217
rect 1233 212 1240 215
rect 1246 217 1253 219
rect 1246 215 1248 217
rect 1250 215 1253 217
rect 1246 212 1253 215
rect 1255 224 1264 226
rect 1255 222 1259 224
rect 1261 222 1264 224
rect 1255 212 1264 222
rect 1222 206 1229 212
rect 1257 206 1264 212
rect 1266 206 1271 226
rect 1273 219 1278 226
rect 1316 223 1321 226
rect 1306 220 1311 223
rect 1273 217 1280 219
rect 1273 215 1276 217
rect 1278 215 1280 217
rect 1273 213 1280 215
rect 1284 217 1291 220
rect 1284 215 1286 217
rect 1288 215 1291 217
rect 1273 206 1278 213
rect 1284 210 1291 215
rect 1284 208 1286 210
rect 1288 208 1291 210
rect 1284 206 1291 208
rect 1293 210 1301 220
rect 1293 208 1296 210
rect 1298 208 1301 210
rect 1293 206 1301 208
rect 1303 218 1311 220
rect 1303 216 1306 218
rect 1308 216 1311 218
rect 1303 213 1311 216
rect 1313 221 1321 223
rect 1313 219 1316 221
rect 1318 219 1321 221
rect 1313 213 1321 219
rect 1323 219 1328 226
rect 1335 223 1341 225
rect 1335 221 1337 223
rect 1339 221 1341 223
rect 1335 219 1341 221
rect 1354 223 1360 225
rect 1401 227 1408 229
rect 1401 225 1404 227
rect 1406 225 1408 227
rect 1354 221 1356 223
rect 1358 221 1360 223
rect 1354 219 1360 221
rect 1323 217 1330 219
rect 1323 215 1326 217
rect 1328 215 1330 217
rect 1323 213 1330 215
rect 1303 206 1308 213
rect 1335 212 1340 219
rect 1356 215 1360 219
rect 1401 219 1408 225
rect 1383 217 1390 219
rect 1383 215 1385 217
rect 1387 215 1390 217
rect 1356 212 1362 215
rect 1335 206 1342 212
rect 1344 210 1352 212
rect 1344 208 1347 210
rect 1349 208 1352 210
rect 1344 206 1352 208
rect 1354 206 1362 212
rect 1364 212 1369 215
rect 1383 213 1390 215
rect 1364 210 1371 212
rect 1364 208 1367 210
rect 1369 208 1371 210
rect 1385 208 1390 213
rect 1392 208 1397 219
rect 1399 217 1408 219
rect 1425 219 1430 226
rect 1423 217 1430 219
rect 1399 208 1410 217
rect 1412 215 1419 217
rect 1412 213 1415 215
rect 1417 213 1419 215
rect 1423 215 1425 217
rect 1427 215 1430 217
rect 1423 213 1430 215
rect 1432 223 1437 226
rect 1432 221 1440 223
rect 1432 219 1435 221
rect 1437 219 1440 221
rect 1432 213 1440 219
rect 1442 220 1447 223
rect 1442 218 1450 220
rect 1442 216 1445 218
rect 1447 216 1450 218
rect 1442 213 1450 216
rect 1412 211 1419 213
rect 1412 208 1417 211
rect 1364 206 1371 208
rect 1445 206 1450 213
rect 1452 210 1460 220
rect 1452 208 1455 210
rect 1457 208 1460 210
rect 1452 206 1460 208
rect 1462 217 1469 220
rect 1475 219 1480 226
rect 1462 215 1465 217
rect 1467 215 1469 217
rect 1462 210 1469 215
rect 1473 217 1480 219
rect 1473 215 1475 217
rect 1477 215 1480 217
rect 1473 213 1480 215
rect 1462 208 1465 210
rect 1467 208 1469 210
rect 1462 206 1469 208
rect 1475 206 1480 213
rect 1482 206 1487 226
rect 1489 224 1498 226
rect 1489 222 1492 224
rect 1494 222 1498 224
rect 1489 212 1498 222
rect 1500 219 1505 226
rect 1515 219 1520 226
rect 1500 217 1507 219
rect 1500 215 1503 217
rect 1505 215 1507 217
rect 1500 212 1507 215
rect 1513 217 1520 219
rect 1513 215 1515 217
rect 1517 215 1520 217
rect 1513 212 1520 215
rect 1522 224 1531 226
rect 1522 222 1526 224
rect 1528 222 1531 224
rect 1522 212 1531 222
rect 1489 206 1496 212
rect 1524 206 1531 212
rect 1533 206 1538 226
rect 1540 219 1545 226
rect 1583 223 1588 226
rect 1573 220 1578 223
rect 1540 217 1547 219
rect 1540 215 1543 217
rect 1545 215 1547 217
rect 1540 213 1547 215
rect 1551 217 1558 220
rect 1551 215 1553 217
rect 1555 215 1558 217
rect 1540 206 1545 213
rect 1551 210 1558 215
rect 1551 208 1553 210
rect 1555 208 1558 210
rect 1551 206 1558 208
rect 1560 210 1568 220
rect 1560 208 1563 210
rect 1565 208 1568 210
rect 1560 206 1568 208
rect 1570 218 1578 220
rect 1570 216 1573 218
rect 1575 216 1578 218
rect 1570 213 1578 216
rect 1580 221 1588 223
rect 1580 219 1583 221
rect 1585 219 1588 221
rect 1580 213 1588 219
rect 1590 219 1595 226
rect 1602 223 1608 225
rect 1602 221 1604 223
rect 1606 221 1608 223
rect 1602 219 1608 221
rect 1621 223 1627 225
rect 1668 227 1675 229
rect 1668 225 1671 227
rect 1673 225 1675 227
rect 1621 221 1623 223
rect 1625 221 1627 223
rect 1621 219 1627 221
rect 1590 217 1597 219
rect 1590 215 1593 217
rect 1595 215 1597 217
rect 1590 213 1597 215
rect 1570 206 1575 213
rect 1602 212 1607 219
rect 1623 215 1627 219
rect 1668 219 1675 225
rect 1650 217 1657 219
rect 1650 215 1652 217
rect 1654 215 1657 217
rect 1623 212 1629 215
rect 1602 206 1609 212
rect 1611 210 1619 212
rect 1611 208 1614 210
rect 1616 208 1619 210
rect 1611 206 1619 208
rect 1621 206 1629 212
rect 1631 212 1636 215
rect 1650 213 1657 215
rect 1631 210 1638 212
rect 1631 208 1634 210
rect 1636 208 1638 210
rect 1652 208 1657 213
rect 1659 208 1664 219
rect 1666 217 1675 219
rect 1692 219 1697 226
rect 1690 217 1697 219
rect 1666 208 1677 217
rect 1679 215 1686 217
rect 1679 213 1682 215
rect 1684 213 1686 215
rect 1690 215 1692 217
rect 1694 215 1697 217
rect 1690 213 1697 215
rect 1699 223 1704 226
rect 1699 221 1707 223
rect 1699 219 1702 221
rect 1704 219 1707 221
rect 1699 213 1707 219
rect 1709 220 1714 223
rect 1709 218 1717 220
rect 1709 216 1712 218
rect 1714 216 1717 218
rect 1709 213 1717 216
rect 1679 211 1686 213
rect 1679 208 1684 211
rect 1631 206 1638 208
rect 1712 206 1717 213
rect 1719 210 1727 220
rect 1719 208 1722 210
rect 1724 208 1727 210
rect 1719 206 1727 208
rect 1729 217 1736 220
rect 1742 219 1747 226
rect 1729 215 1732 217
rect 1734 215 1736 217
rect 1729 210 1736 215
rect 1740 217 1747 219
rect 1740 215 1742 217
rect 1744 215 1747 217
rect 1740 213 1747 215
rect 1729 208 1732 210
rect 1734 208 1736 210
rect 1729 206 1736 208
rect 1742 206 1747 213
rect 1749 206 1754 226
rect 1756 224 1765 226
rect 1756 222 1759 224
rect 1761 222 1765 224
rect 1756 212 1765 222
rect 1767 219 1772 226
rect 1782 219 1787 226
rect 1767 217 1774 219
rect 1767 215 1770 217
rect 1772 215 1774 217
rect 1767 212 1774 215
rect 1780 217 1787 219
rect 1780 215 1782 217
rect 1784 215 1787 217
rect 1780 212 1787 215
rect 1789 224 1798 226
rect 1789 222 1793 224
rect 1795 222 1798 224
rect 1789 212 1798 222
rect 1756 206 1763 212
rect 1791 206 1798 212
rect 1800 206 1805 226
rect 1807 219 1812 226
rect 1850 223 1855 226
rect 1840 220 1845 223
rect 1807 217 1814 219
rect 1807 215 1810 217
rect 1812 215 1814 217
rect 1807 213 1814 215
rect 1818 217 1825 220
rect 1818 215 1820 217
rect 1822 215 1825 217
rect 1807 206 1812 213
rect 1818 210 1825 215
rect 1818 208 1820 210
rect 1822 208 1825 210
rect 1818 206 1825 208
rect 1827 210 1835 220
rect 1827 208 1830 210
rect 1832 208 1835 210
rect 1827 206 1835 208
rect 1837 218 1845 220
rect 1837 216 1840 218
rect 1842 216 1845 218
rect 1837 213 1845 216
rect 1847 221 1855 223
rect 1847 219 1850 221
rect 1852 219 1855 221
rect 1847 213 1855 219
rect 1857 219 1862 226
rect 1869 223 1875 225
rect 1869 221 1871 223
rect 1873 221 1875 223
rect 1869 219 1875 221
rect 1888 223 1894 225
rect 1888 221 1890 223
rect 1892 221 1894 223
rect 1888 219 1894 221
rect 1966 227 1972 229
rect 1966 225 1968 227
rect 1970 225 1972 227
rect 1966 223 1972 225
rect 1950 220 1955 223
rect 1857 217 1864 219
rect 1857 215 1860 217
rect 1862 215 1864 217
rect 1857 213 1864 215
rect 1837 206 1842 213
rect 1869 212 1874 219
rect 1890 215 1894 219
rect 1926 218 1935 220
rect 1926 216 1928 218
rect 1930 216 1935 218
rect 1926 215 1935 216
rect 1890 212 1896 215
rect 1869 206 1876 212
rect 1878 210 1886 212
rect 1878 208 1881 210
rect 1883 208 1886 210
rect 1878 206 1886 208
rect 1888 206 1896 212
rect 1898 212 1903 215
rect 1914 212 1919 215
rect 1898 210 1905 212
rect 1898 208 1901 210
rect 1903 208 1905 210
rect 1898 206 1905 208
rect 1912 210 1919 212
rect 1912 208 1914 210
rect 1916 208 1919 210
rect 1912 206 1919 208
rect 1921 211 1935 215
rect 1937 215 1945 220
rect 1937 213 1940 215
rect 1942 213 1945 215
rect 1937 211 1945 213
rect 1947 217 1955 220
rect 1947 215 1950 217
rect 1952 215 1955 217
rect 1947 211 1955 215
rect 1957 211 1962 223
rect 1964 211 1972 223
rect 1978 219 1983 226
rect 1976 217 1983 219
rect 1976 215 1978 217
rect 1980 215 1983 217
rect 1976 213 1983 215
rect 1985 223 1990 226
rect 1985 221 1993 223
rect 1985 219 1988 221
rect 1990 219 1993 221
rect 1985 213 1993 219
rect 1995 220 2000 223
rect 1995 218 2003 220
rect 1995 216 1998 218
rect 2000 216 2003 218
rect 1995 213 2003 216
rect 1921 206 1926 211
rect 1998 206 2003 213
rect 2005 210 2013 220
rect 2005 208 2008 210
rect 2010 208 2013 210
rect 2005 206 2013 208
rect 2015 217 2022 220
rect 2028 219 2033 226
rect 2015 215 2018 217
rect 2020 215 2022 217
rect 2015 210 2022 215
rect 2026 217 2033 219
rect 2026 215 2028 217
rect 2030 215 2033 217
rect 2026 213 2033 215
rect 2015 208 2018 210
rect 2020 208 2022 210
rect 2015 206 2022 208
rect 2028 206 2033 213
rect 2035 206 2040 226
rect 2042 224 2051 226
rect 2042 222 2045 224
rect 2047 222 2051 224
rect 2042 212 2051 222
rect 2053 219 2058 226
rect 2068 219 2073 226
rect 2053 217 2060 219
rect 2053 215 2056 217
rect 2058 215 2060 217
rect 2053 212 2060 215
rect 2066 217 2073 219
rect 2066 215 2068 217
rect 2070 215 2073 217
rect 2066 212 2073 215
rect 2075 224 2084 226
rect 2075 222 2079 224
rect 2081 222 2084 224
rect 2075 212 2084 222
rect 2042 206 2049 212
rect 2077 206 2084 212
rect 2086 206 2091 226
rect 2093 219 2098 226
rect 2136 223 2141 226
rect 2126 220 2131 223
rect 2093 217 2100 219
rect 2093 215 2096 217
rect 2098 215 2100 217
rect 2093 213 2100 215
rect 2104 217 2111 220
rect 2104 215 2106 217
rect 2108 215 2111 217
rect 2093 206 2098 213
rect 2104 210 2111 215
rect 2104 208 2106 210
rect 2108 208 2111 210
rect 2104 206 2111 208
rect 2113 210 2121 220
rect 2113 208 2116 210
rect 2118 208 2121 210
rect 2113 206 2121 208
rect 2123 218 2131 220
rect 2123 216 2126 218
rect 2128 216 2131 218
rect 2123 213 2131 216
rect 2133 221 2141 223
rect 2133 219 2136 221
rect 2138 219 2141 221
rect 2133 213 2141 219
rect 2143 219 2148 226
rect 2155 223 2161 225
rect 2155 221 2157 223
rect 2159 221 2161 223
rect 2155 219 2161 221
rect 2174 223 2180 225
rect 2174 221 2176 223
rect 2178 221 2180 223
rect 2174 219 2180 221
rect 2143 217 2150 219
rect 2143 215 2146 217
rect 2148 215 2150 217
rect 2143 213 2150 215
rect 2123 206 2128 213
rect 2155 212 2160 219
rect 2176 215 2180 219
rect 2210 218 2216 220
rect 2199 216 2206 218
rect 2176 212 2182 215
rect 2155 206 2162 212
rect 2164 210 2172 212
rect 2164 208 2167 210
rect 2169 208 2172 210
rect 2164 206 2172 208
rect 2174 206 2182 212
rect 2184 212 2189 215
rect 2199 214 2201 216
rect 2203 214 2206 216
rect 2199 212 2206 214
rect 2208 216 2216 218
rect 2208 214 2211 216
rect 2213 214 2216 216
rect 2208 212 2216 214
rect 2218 212 2223 220
rect 2225 218 2233 220
rect 2225 216 2228 218
rect 2230 216 2233 218
rect 2225 212 2233 216
rect 2235 212 2240 220
rect 2242 218 2250 220
rect 2242 216 2245 218
rect 2247 216 2250 218
rect 2242 212 2250 216
rect 2184 210 2191 212
rect 2184 208 2187 210
rect 2189 208 2191 210
rect 2184 206 2191 208
rect 2245 211 2250 212
rect 2252 217 2257 220
rect 2278 218 2284 220
rect 2252 215 2259 217
rect 2252 213 2255 215
rect 2257 213 2259 215
rect 2252 211 2259 213
rect 2267 216 2274 218
rect 2267 214 2269 216
rect 2271 214 2274 216
rect 2267 212 2274 214
rect 2276 216 2284 218
rect 2276 214 2279 216
rect 2281 214 2284 216
rect 2276 212 2284 214
rect 2286 212 2291 220
rect 2293 218 2301 220
rect 2293 216 2296 218
rect 2298 216 2301 218
rect 2293 212 2301 216
rect 2303 212 2308 220
rect 2310 218 2318 220
rect 2310 216 2313 218
rect 2315 216 2318 218
rect 2310 212 2318 216
rect 2313 211 2318 212
rect 2320 217 2325 220
rect 2320 215 2327 217
rect 2320 213 2323 215
rect 2325 213 2327 215
rect 2320 211 2327 213
rect 10 107 15 112
rect 8 105 15 107
rect 8 103 10 105
rect 12 103 15 105
rect 8 101 15 103
rect 17 101 22 112
rect 24 103 35 112
rect 37 109 42 112
rect 37 107 44 109
rect 50 107 55 112
rect 37 105 40 107
rect 42 105 44 107
rect 37 103 44 105
rect 48 105 55 107
rect 48 103 50 105
rect 52 103 55 105
rect 24 101 33 103
rect 26 95 33 101
rect 48 101 55 103
rect 57 101 62 112
rect 64 103 75 112
rect 77 109 82 112
rect 77 107 84 109
rect 110 107 115 114
rect 77 105 80 107
rect 82 105 84 107
rect 77 103 84 105
rect 88 105 95 107
rect 88 103 90 105
rect 92 103 95 105
rect 64 101 73 103
rect 26 93 29 95
rect 31 93 33 95
rect 26 91 33 93
rect 66 95 73 101
rect 88 101 95 103
rect 66 93 69 95
rect 71 93 73 95
rect 66 91 73 93
rect 90 94 95 101
rect 97 101 105 107
rect 97 99 100 101
rect 102 99 105 101
rect 97 97 105 99
rect 107 104 115 107
rect 107 102 110 104
rect 112 102 115 104
rect 107 100 115 102
rect 117 112 125 114
rect 117 110 120 112
rect 122 110 125 112
rect 117 100 125 110
rect 127 112 134 114
rect 127 110 130 112
rect 132 110 134 112
rect 127 105 134 110
rect 140 107 145 114
rect 127 103 130 105
rect 132 103 134 105
rect 127 100 134 103
rect 138 105 145 107
rect 138 103 140 105
rect 142 103 145 105
rect 138 101 145 103
rect 107 97 112 100
rect 97 94 102 97
rect 140 94 145 101
rect 147 94 152 114
rect 154 108 161 114
rect 189 108 196 114
rect 154 98 163 108
rect 154 96 157 98
rect 159 96 163 98
rect 154 94 163 96
rect 165 105 172 108
rect 165 103 168 105
rect 170 103 172 105
rect 165 101 172 103
rect 178 105 185 108
rect 178 103 180 105
rect 182 103 185 105
rect 178 101 185 103
rect 165 94 170 101
rect 180 94 185 101
rect 187 98 196 108
rect 187 96 191 98
rect 193 96 196 98
rect 187 94 196 96
rect 198 94 203 114
rect 205 107 210 114
rect 216 112 223 114
rect 216 110 218 112
rect 220 110 223 112
rect 205 105 212 107
rect 205 103 208 105
rect 210 103 212 105
rect 205 101 212 103
rect 216 105 223 110
rect 216 103 218 105
rect 220 103 223 105
rect 205 94 210 101
rect 216 100 223 103
rect 225 112 233 114
rect 225 110 228 112
rect 230 110 233 112
rect 225 100 233 110
rect 235 107 240 114
rect 267 108 274 114
rect 276 112 284 114
rect 276 110 279 112
rect 281 110 284 112
rect 276 108 284 110
rect 286 108 294 114
rect 235 104 243 107
rect 235 102 238 104
rect 240 102 243 104
rect 235 100 243 102
rect 238 97 243 100
rect 245 101 253 107
rect 245 99 248 101
rect 250 99 253 101
rect 245 97 253 99
rect 248 94 253 97
rect 255 105 262 107
rect 255 103 258 105
rect 260 103 262 105
rect 255 101 262 103
rect 267 101 272 108
rect 288 105 294 108
rect 296 112 303 114
rect 296 110 299 112
rect 301 110 303 112
rect 296 108 303 110
rect 296 105 301 108
rect 317 107 322 112
rect 315 105 322 107
rect 288 101 292 105
rect 255 94 260 101
rect 267 99 273 101
rect 267 97 269 99
rect 271 97 273 99
rect 267 95 273 97
rect 286 99 292 101
rect 315 103 317 105
rect 319 103 322 105
rect 315 101 322 103
rect 324 101 329 112
rect 331 103 342 112
rect 344 109 349 112
rect 344 107 351 109
rect 377 107 382 114
rect 344 105 347 107
rect 349 105 351 107
rect 344 103 351 105
rect 355 105 362 107
rect 355 103 357 105
rect 359 103 362 105
rect 331 101 340 103
rect 286 97 288 99
rect 290 97 292 99
rect 286 95 292 97
rect 333 95 340 101
rect 355 101 362 103
rect 333 93 336 95
rect 338 93 340 95
rect 333 91 340 93
rect 357 94 362 101
rect 364 101 372 107
rect 364 99 367 101
rect 369 99 372 101
rect 364 97 372 99
rect 374 104 382 107
rect 374 102 377 104
rect 379 102 382 104
rect 374 100 382 102
rect 384 112 392 114
rect 384 110 387 112
rect 389 110 392 112
rect 384 100 392 110
rect 394 112 401 114
rect 394 110 397 112
rect 399 110 401 112
rect 394 105 401 110
rect 407 107 412 114
rect 394 103 397 105
rect 399 103 401 105
rect 394 100 401 103
rect 405 105 412 107
rect 405 103 407 105
rect 409 103 412 105
rect 405 101 412 103
rect 374 97 379 100
rect 364 94 369 97
rect 407 94 412 101
rect 414 94 419 114
rect 421 108 428 114
rect 456 108 463 114
rect 421 98 430 108
rect 421 96 424 98
rect 426 96 430 98
rect 421 94 430 96
rect 432 105 439 108
rect 432 103 435 105
rect 437 103 439 105
rect 432 101 439 103
rect 445 105 452 108
rect 445 103 447 105
rect 449 103 452 105
rect 445 101 452 103
rect 432 94 437 101
rect 447 94 452 101
rect 454 98 463 108
rect 454 96 458 98
rect 460 96 463 98
rect 454 94 463 96
rect 465 94 470 114
rect 472 107 477 114
rect 483 112 490 114
rect 483 110 485 112
rect 487 110 490 112
rect 472 105 479 107
rect 472 103 475 105
rect 477 103 479 105
rect 472 101 479 103
rect 483 105 490 110
rect 483 103 485 105
rect 487 103 490 105
rect 472 94 477 101
rect 483 100 490 103
rect 492 112 500 114
rect 492 110 495 112
rect 497 110 500 112
rect 492 100 500 110
rect 502 107 507 114
rect 534 108 541 114
rect 543 112 551 114
rect 543 110 546 112
rect 548 110 551 112
rect 543 108 551 110
rect 553 108 561 114
rect 502 104 510 107
rect 502 102 505 104
rect 507 102 510 104
rect 502 100 510 102
rect 505 97 510 100
rect 512 101 520 107
rect 512 99 515 101
rect 517 99 520 101
rect 512 97 520 99
rect 515 94 520 97
rect 522 105 529 107
rect 522 103 525 105
rect 527 103 529 105
rect 522 101 529 103
rect 534 101 539 108
rect 555 105 561 108
rect 563 112 570 114
rect 563 110 566 112
rect 568 110 570 112
rect 563 108 570 110
rect 563 105 568 108
rect 584 107 589 112
rect 582 105 589 107
rect 555 101 559 105
rect 522 94 527 101
rect 534 99 540 101
rect 534 97 536 99
rect 538 97 540 99
rect 534 95 540 97
rect 553 99 559 101
rect 582 103 584 105
rect 586 103 589 105
rect 582 101 589 103
rect 591 101 596 112
rect 598 103 609 112
rect 611 109 616 112
rect 611 107 618 109
rect 644 107 649 114
rect 611 105 614 107
rect 616 105 618 107
rect 611 103 618 105
rect 622 105 629 107
rect 622 103 624 105
rect 626 103 629 105
rect 598 101 607 103
rect 553 97 555 99
rect 557 97 559 99
rect 553 95 559 97
rect 600 95 607 101
rect 622 101 629 103
rect 600 93 603 95
rect 605 93 607 95
rect 600 91 607 93
rect 624 94 629 101
rect 631 101 639 107
rect 631 99 634 101
rect 636 99 639 101
rect 631 97 639 99
rect 641 104 649 107
rect 641 102 644 104
rect 646 102 649 104
rect 641 100 649 102
rect 651 112 659 114
rect 651 110 654 112
rect 656 110 659 112
rect 651 100 659 110
rect 661 112 668 114
rect 661 110 664 112
rect 666 110 668 112
rect 661 105 668 110
rect 674 107 679 114
rect 661 103 664 105
rect 666 103 668 105
rect 661 100 668 103
rect 672 105 679 107
rect 672 103 674 105
rect 676 103 679 105
rect 672 101 679 103
rect 641 97 646 100
rect 631 94 636 97
rect 674 94 679 101
rect 681 94 686 114
rect 688 108 695 114
rect 723 108 730 114
rect 688 98 697 108
rect 688 96 691 98
rect 693 96 697 98
rect 688 94 697 96
rect 699 105 706 108
rect 699 103 702 105
rect 704 103 706 105
rect 699 101 706 103
rect 712 105 719 108
rect 712 103 714 105
rect 716 103 719 105
rect 712 101 719 103
rect 699 94 704 101
rect 714 94 719 101
rect 721 98 730 108
rect 721 96 725 98
rect 727 96 730 98
rect 721 94 730 96
rect 732 94 737 114
rect 739 107 744 114
rect 750 112 757 114
rect 750 110 752 112
rect 754 110 757 112
rect 739 105 746 107
rect 739 103 742 105
rect 744 103 746 105
rect 739 101 746 103
rect 750 105 757 110
rect 750 103 752 105
rect 754 103 757 105
rect 739 94 744 101
rect 750 100 757 103
rect 759 112 767 114
rect 759 110 762 112
rect 764 110 767 112
rect 759 100 767 110
rect 769 107 774 114
rect 801 108 808 114
rect 810 112 818 114
rect 810 110 813 112
rect 815 110 818 112
rect 810 108 818 110
rect 820 108 828 114
rect 769 104 777 107
rect 769 102 772 104
rect 774 102 777 104
rect 769 100 777 102
rect 772 97 777 100
rect 779 101 787 107
rect 779 99 782 101
rect 784 99 787 101
rect 779 97 787 99
rect 782 94 787 97
rect 789 105 796 107
rect 789 103 792 105
rect 794 103 796 105
rect 789 101 796 103
rect 801 101 806 108
rect 822 105 828 108
rect 830 112 837 114
rect 830 110 833 112
rect 835 110 837 112
rect 830 108 837 110
rect 830 105 835 108
rect 851 107 856 112
rect 849 105 856 107
rect 822 101 826 105
rect 789 94 794 101
rect 801 99 807 101
rect 801 97 803 99
rect 805 97 807 99
rect 801 95 807 97
rect 820 99 826 101
rect 849 103 851 105
rect 853 103 856 105
rect 849 101 856 103
rect 858 101 863 112
rect 865 103 876 112
rect 878 109 883 112
rect 878 107 885 109
rect 911 107 916 114
rect 878 105 881 107
rect 883 105 885 107
rect 878 103 885 105
rect 889 105 896 107
rect 889 103 891 105
rect 893 103 896 105
rect 865 101 874 103
rect 820 97 822 99
rect 824 97 826 99
rect 820 95 826 97
rect 867 95 874 101
rect 889 101 896 103
rect 867 93 870 95
rect 872 93 874 95
rect 867 91 874 93
rect 891 94 896 101
rect 898 101 906 107
rect 898 99 901 101
rect 903 99 906 101
rect 898 97 906 99
rect 908 104 916 107
rect 908 102 911 104
rect 913 102 916 104
rect 908 100 916 102
rect 918 112 926 114
rect 918 110 921 112
rect 923 110 926 112
rect 918 100 926 110
rect 928 112 935 114
rect 928 110 931 112
rect 933 110 935 112
rect 928 105 935 110
rect 941 107 946 114
rect 928 103 931 105
rect 933 103 935 105
rect 928 100 935 103
rect 939 105 946 107
rect 939 103 941 105
rect 943 103 946 105
rect 939 101 946 103
rect 908 97 913 100
rect 898 94 903 97
rect 941 94 946 101
rect 948 94 953 114
rect 955 108 962 114
rect 990 108 997 114
rect 955 98 964 108
rect 955 96 958 98
rect 960 96 964 98
rect 955 94 964 96
rect 966 105 973 108
rect 966 103 969 105
rect 971 103 973 105
rect 966 101 973 103
rect 979 105 986 108
rect 979 103 981 105
rect 983 103 986 105
rect 979 101 986 103
rect 966 94 971 101
rect 981 94 986 101
rect 988 98 997 108
rect 988 96 992 98
rect 994 96 997 98
rect 988 94 997 96
rect 999 94 1004 114
rect 1006 107 1011 114
rect 1017 112 1024 114
rect 1017 110 1019 112
rect 1021 110 1024 112
rect 1006 105 1013 107
rect 1006 103 1009 105
rect 1011 103 1013 105
rect 1006 101 1013 103
rect 1017 105 1024 110
rect 1017 103 1019 105
rect 1021 103 1024 105
rect 1006 94 1011 101
rect 1017 100 1024 103
rect 1026 112 1034 114
rect 1026 110 1029 112
rect 1031 110 1034 112
rect 1026 100 1034 110
rect 1036 107 1041 114
rect 1068 108 1075 114
rect 1077 112 1085 114
rect 1077 110 1080 112
rect 1082 110 1085 112
rect 1077 108 1085 110
rect 1087 108 1095 114
rect 1036 104 1044 107
rect 1036 102 1039 104
rect 1041 102 1044 104
rect 1036 100 1044 102
rect 1039 97 1044 100
rect 1046 101 1054 107
rect 1046 99 1049 101
rect 1051 99 1054 101
rect 1046 97 1054 99
rect 1049 94 1054 97
rect 1056 105 1063 107
rect 1056 103 1059 105
rect 1061 103 1063 105
rect 1056 101 1063 103
rect 1068 101 1073 108
rect 1089 105 1095 108
rect 1097 112 1104 114
rect 1097 110 1100 112
rect 1102 110 1104 112
rect 1097 108 1104 110
rect 1097 105 1102 108
rect 1118 107 1123 112
rect 1116 105 1123 107
rect 1089 101 1093 105
rect 1056 94 1061 101
rect 1068 99 1074 101
rect 1068 97 1070 99
rect 1072 97 1074 99
rect 1068 95 1074 97
rect 1087 99 1093 101
rect 1116 103 1118 105
rect 1120 103 1123 105
rect 1116 101 1123 103
rect 1125 101 1130 112
rect 1132 103 1143 112
rect 1145 109 1150 112
rect 1145 107 1152 109
rect 1178 107 1183 114
rect 1145 105 1148 107
rect 1150 105 1152 107
rect 1145 103 1152 105
rect 1156 105 1163 107
rect 1156 103 1158 105
rect 1160 103 1163 105
rect 1132 101 1141 103
rect 1087 97 1089 99
rect 1091 97 1093 99
rect 1087 95 1093 97
rect 1134 95 1141 101
rect 1156 101 1163 103
rect 1134 93 1137 95
rect 1139 93 1141 95
rect 1134 91 1141 93
rect 1158 94 1163 101
rect 1165 101 1173 107
rect 1165 99 1168 101
rect 1170 99 1173 101
rect 1165 97 1173 99
rect 1175 104 1183 107
rect 1175 102 1178 104
rect 1180 102 1183 104
rect 1175 100 1183 102
rect 1185 112 1193 114
rect 1185 110 1188 112
rect 1190 110 1193 112
rect 1185 100 1193 110
rect 1195 112 1202 114
rect 1195 110 1198 112
rect 1200 110 1202 112
rect 1195 105 1202 110
rect 1208 107 1213 114
rect 1195 103 1198 105
rect 1200 103 1202 105
rect 1195 100 1202 103
rect 1206 105 1213 107
rect 1206 103 1208 105
rect 1210 103 1213 105
rect 1206 101 1213 103
rect 1175 97 1180 100
rect 1165 94 1170 97
rect 1208 94 1213 101
rect 1215 94 1220 114
rect 1222 108 1229 114
rect 1257 108 1264 114
rect 1222 98 1231 108
rect 1222 96 1225 98
rect 1227 96 1231 98
rect 1222 94 1231 96
rect 1233 105 1240 108
rect 1233 103 1236 105
rect 1238 103 1240 105
rect 1233 101 1240 103
rect 1246 105 1253 108
rect 1246 103 1248 105
rect 1250 103 1253 105
rect 1246 101 1253 103
rect 1233 94 1238 101
rect 1248 94 1253 101
rect 1255 98 1264 108
rect 1255 96 1259 98
rect 1261 96 1264 98
rect 1255 94 1264 96
rect 1266 94 1271 114
rect 1273 107 1278 114
rect 1284 112 1291 114
rect 1284 110 1286 112
rect 1288 110 1291 112
rect 1273 105 1280 107
rect 1273 103 1276 105
rect 1278 103 1280 105
rect 1273 101 1280 103
rect 1284 105 1291 110
rect 1284 103 1286 105
rect 1288 103 1291 105
rect 1273 94 1278 101
rect 1284 100 1291 103
rect 1293 112 1301 114
rect 1293 110 1296 112
rect 1298 110 1301 112
rect 1293 100 1301 110
rect 1303 107 1308 114
rect 1335 108 1342 114
rect 1344 112 1352 114
rect 1344 110 1347 112
rect 1349 110 1352 112
rect 1344 108 1352 110
rect 1354 108 1362 114
rect 1303 104 1311 107
rect 1303 102 1306 104
rect 1308 102 1311 104
rect 1303 100 1311 102
rect 1306 97 1311 100
rect 1313 101 1321 107
rect 1313 99 1316 101
rect 1318 99 1321 101
rect 1313 97 1321 99
rect 1316 94 1321 97
rect 1323 105 1330 107
rect 1323 103 1326 105
rect 1328 103 1330 105
rect 1323 101 1330 103
rect 1335 101 1340 108
rect 1356 105 1362 108
rect 1364 112 1371 114
rect 1364 110 1367 112
rect 1369 110 1371 112
rect 1364 108 1371 110
rect 1364 105 1369 108
rect 1385 107 1390 112
rect 1383 105 1390 107
rect 1356 101 1360 105
rect 1323 94 1328 101
rect 1335 99 1341 101
rect 1335 97 1337 99
rect 1339 97 1341 99
rect 1335 95 1341 97
rect 1354 99 1360 101
rect 1383 103 1385 105
rect 1387 103 1390 105
rect 1383 101 1390 103
rect 1392 101 1397 112
rect 1399 103 1410 112
rect 1412 109 1417 112
rect 1412 107 1419 109
rect 1445 107 1450 114
rect 1412 105 1415 107
rect 1417 105 1419 107
rect 1412 103 1419 105
rect 1423 105 1430 107
rect 1423 103 1425 105
rect 1427 103 1430 105
rect 1399 101 1408 103
rect 1354 97 1356 99
rect 1358 97 1360 99
rect 1354 95 1360 97
rect 1401 95 1408 101
rect 1423 101 1430 103
rect 1401 93 1404 95
rect 1406 93 1408 95
rect 1401 91 1408 93
rect 1425 94 1430 101
rect 1432 101 1440 107
rect 1432 99 1435 101
rect 1437 99 1440 101
rect 1432 97 1440 99
rect 1442 104 1450 107
rect 1442 102 1445 104
rect 1447 102 1450 104
rect 1442 100 1450 102
rect 1452 112 1460 114
rect 1452 110 1455 112
rect 1457 110 1460 112
rect 1452 100 1460 110
rect 1462 112 1469 114
rect 1462 110 1465 112
rect 1467 110 1469 112
rect 1462 105 1469 110
rect 1475 107 1480 114
rect 1462 103 1465 105
rect 1467 103 1469 105
rect 1462 100 1469 103
rect 1473 105 1480 107
rect 1473 103 1475 105
rect 1477 103 1480 105
rect 1473 101 1480 103
rect 1442 97 1447 100
rect 1432 94 1437 97
rect 1475 94 1480 101
rect 1482 94 1487 114
rect 1489 108 1496 114
rect 1524 108 1531 114
rect 1489 98 1498 108
rect 1489 96 1492 98
rect 1494 96 1498 98
rect 1489 94 1498 96
rect 1500 105 1507 108
rect 1500 103 1503 105
rect 1505 103 1507 105
rect 1500 101 1507 103
rect 1513 105 1520 108
rect 1513 103 1515 105
rect 1517 103 1520 105
rect 1513 101 1520 103
rect 1500 94 1505 101
rect 1515 94 1520 101
rect 1522 98 1531 108
rect 1522 96 1526 98
rect 1528 96 1531 98
rect 1522 94 1531 96
rect 1533 94 1538 114
rect 1540 107 1545 114
rect 1551 112 1558 114
rect 1551 110 1553 112
rect 1555 110 1558 112
rect 1540 105 1547 107
rect 1540 103 1543 105
rect 1545 103 1547 105
rect 1540 101 1547 103
rect 1551 105 1558 110
rect 1551 103 1553 105
rect 1555 103 1558 105
rect 1540 94 1545 101
rect 1551 100 1558 103
rect 1560 112 1568 114
rect 1560 110 1563 112
rect 1565 110 1568 112
rect 1560 100 1568 110
rect 1570 107 1575 114
rect 1602 108 1609 114
rect 1611 112 1619 114
rect 1611 110 1614 112
rect 1616 110 1619 112
rect 1611 108 1619 110
rect 1621 108 1629 114
rect 1570 104 1578 107
rect 1570 102 1573 104
rect 1575 102 1578 104
rect 1570 100 1578 102
rect 1573 97 1578 100
rect 1580 101 1588 107
rect 1580 99 1583 101
rect 1585 99 1588 101
rect 1580 97 1588 99
rect 1583 94 1588 97
rect 1590 105 1597 107
rect 1590 103 1593 105
rect 1595 103 1597 105
rect 1590 101 1597 103
rect 1602 101 1607 108
rect 1623 105 1629 108
rect 1631 112 1638 114
rect 1631 110 1634 112
rect 1636 110 1638 112
rect 1631 108 1638 110
rect 1631 105 1636 108
rect 1652 107 1657 112
rect 1650 105 1657 107
rect 1623 101 1627 105
rect 1590 94 1595 101
rect 1602 99 1608 101
rect 1602 97 1604 99
rect 1606 97 1608 99
rect 1602 95 1608 97
rect 1621 99 1627 101
rect 1650 103 1652 105
rect 1654 103 1657 105
rect 1650 101 1657 103
rect 1659 101 1664 112
rect 1666 103 1677 112
rect 1679 109 1684 112
rect 1679 107 1686 109
rect 1712 107 1717 114
rect 1679 105 1682 107
rect 1684 105 1686 107
rect 1679 103 1686 105
rect 1690 105 1697 107
rect 1690 103 1692 105
rect 1694 103 1697 105
rect 1666 101 1675 103
rect 1621 97 1623 99
rect 1625 97 1627 99
rect 1621 95 1627 97
rect 1668 95 1675 101
rect 1690 101 1697 103
rect 1668 93 1671 95
rect 1673 93 1675 95
rect 1668 91 1675 93
rect 1692 94 1697 101
rect 1699 101 1707 107
rect 1699 99 1702 101
rect 1704 99 1707 101
rect 1699 97 1707 99
rect 1709 104 1717 107
rect 1709 102 1712 104
rect 1714 102 1717 104
rect 1709 100 1717 102
rect 1719 112 1727 114
rect 1719 110 1722 112
rect 1724 110 1727 112
rect 1719 100 1727 110
rect 1729 112 1736 114
rect 1729 110 1732 112
rect 1734 110 1736 112
rect 1729 105 1736 110
rect 1742 107 1747 114
rect 1729 103 1732 105
rect 1734 103 1736 105
rect 1729 100 1736 103
rect 1740 105 1747 107
rect 1740 103 1742 105
rect 1744 103 1747 105
rect 1740 101 1747 103
rect 1709 97 1714 100
rect 1699 94 1704 97
rect 1742 94 1747 101
rect 1749 94 1754 114
rect 1756 108 1763 114
rect 1791 108 1798 114
rect 1756 98 1765 108
rect 1756 96 1759 98
rect 1761 96 1765 98
rect 1756 94 1765 96
rect 1767 105 1774 108
rect 1767 103 1770 105
rect 1772 103 1774 105
rect 1767 101 1774 103
rect 1780 105 1787 108
rect 1780 103 1782 105
rect 1784 103 1787 105
rect 1780 101 1787 103
rect 1767 94 1772 101
rect 1782 94 1787 101
rect 1789 98 1798 108
rect 1789 96 1793 98
rect 1795 96 1798 98
rect 1789 94 1798 96
rect 1800 94 1805 114
rect 1807 107 1812 114
rect 1818 112 1825 114
rect 1818 110 1820 112
rect 1822 110 1825 112
rect 1807 105 1814 107
rect 1807 103 1810 105
rect 1812 103 1814 105
rect 1807 101 1814 103
rect 1818 105 1825 110
rect 1818 103 1820 105
rect 1822 103 1825 105
rect 1807 94 1812 101
rect 1818 100 1825 103
rect 1827 112 1835 114
rect 1827 110 1830 112
rect 1832 110 1835 112
rect 1827 100 1835 110
rect 1837 107 1842 114
rect 1869 108 1876 114
rect 1878 112 1886 114
rect 1878 110 1881 112
rect 1883 110 1886 112
rect 1878 108 1886 110
rect 1888 108 1896 114
rect 1837 104 1845 107
rect 1837 102 1840 104
rect 1842 102 1845 104
rect 1837 100 1845 102
rect 1840 97 1845 100
rect 1847 101 1855 107
rect 1847 99 1850 101
rect 1852 99 1855 101
rect 1847 97 1855 99
rect 1850 94 1855 97
rect 1857 105 1864 107
rect 1857 103 1860 105
rect 1862 103 1864 105
rect 1857 101 1864 103
rect 1869 101 1874 108
rect 1890 105 1896 108
rect 1898 112 1905 114
rect 1898 110 1901 112
rect 1903 110 1905 112
rect 1898 108 1905 110
rect 1912 112 1919 114
rect 1912 110 1914 112
rect 1916 110 1919 112
rect 1912 108 1919 110
rect 1898 105 1903 108
rect 1914 105 1919 108
rect 1921 109 1926 114
rect 1921 105 1935 109
rect 1890 101 1894 105
rect 1857 94 1862 101
rect 1869 99 1875 101
rect 1869 97 1871 99
rect 1873 97 1875 99
rect 1869 95 1875 97
rect 1888 99 1894 101
rect 1926 104 1935 105
rect 1926 102 1928 104
rect 1930 102 1935 104
rect 1926 100 1935 102
rect 1937 107 1945 109
rect 1937 105 1940 107
rect 1942 105 1945 107
rect 1937 100 1945 105
rect 1947 105 1955 109
rect 1947 103 1950 105
rect 1952 103 1955 105
rect 1947 100 1955 103
rect 1888 97 1890 99
rect 1892 97 1894 99
rect 1888 95 1894 97
rect 1950 97 1955 100
rect 1957 97 1962 109
rect 1964 97 1972 109
rect 1998 107 2003 114
rect 1976 105 1983 107
rect 1976 103 1978 105
rect 1980 103 1983 105
rect 1976 101 1983 103
rect 1966 95 1972 97
rect 1966 93 1968 95
rect 1970 93 1972 95
rect 1978 94 1983 101
rect 1985 101 1993 107
rect 1985 99 1988 101
rect 1990 99 1993 101
rect 1985 97 1993 99
rect 1995 104 2003 107
rect 1995 102 1998 104
rect 2000 102 2003 104
rect 1995 100 2003 102
rect 2005 112 2013 114
rect 2005 110 2008 112
rect 2010 110 2013 112
rect 2005 100 2013 110
rect 2015 112 2022 114
rect 2015 110 2018 112
rect 2020 110 2022 112
rect 2015 105 2022 110
rect 2028 107 2033 114
rect 2015 103 2018 105
rect 2020 103 2022 105
rect 2015 100 2022 103
rect 2026 105 2033 107
rect 2026 103 2028 105
rect 2030 103 2033 105
rect 2026 101 2033 103
rect 1995 97 2000 100
rect 1985 94 1990 97
rect 1966 91 1972 93
rect 2028 94 2033 101
rect 2035 94 2040 114
rect 2042 108 2049 114
rect 2077 108 2084 114
rect 2042 98 2051 108
rect 2042 96 2045 98
rect 2047 96 2051 98
rect 2042 94 2051 96
rect 2053 105 2060 108
rect 2053 103 2056 105
rect 2058 103 2060 105
rect 2053 101 2060 103
rect 2066 105 2073 108
rect 2066 103 2068 105
rect 2070 103 2073 105
rect 2066 101 2073 103
rect 2053 94 2058 101
rect 2068 94 2073 101
rect 2075 98 2084 108
rect 2075 96 2079 98
rect 2081 96 2084 98
rect 2075 94 2084 96
rect 2086 94 2091 114
rect 2093 107 2098 114
rect 2104 112 2111 114
rect 2104 110 2106 112
rect 2108 110 2111 112
rect 2093 105 2100 107
rect 2093 103 2096 105
rect 2098 103 2100 105
rect 2093 101 2100 103
rect 2104 105 2111 110
rect 2104 103 2106 105
rect 2108 103 2111 105
rect 2093 94 2098 101
rect 2104 100 2111 103
rect 2113 112 2121 114
rect 2113 110 2116 112
rect 2118 110 2121 112
rect 2113 100 2121 110
rect 2123 107 2128 114
rect 2155 108 2162 114
rect 2164 112 2172 114
rect 2164 110 2167 112
rect 2169 110 2172 112
rect 2164 108 2172 110
rect 2174 108 2182 114
rect 2123 104 2131 107
rect 2123 102 2126 104
rect 2128 102 2131 104
rect 2123 100 2131 102
rect 2126 97 2131 100
rect 2133 101 2141 107
rect 2133 99 2136 101
rect 2138 99 2141 101
rect 2133 97 2141 99
rect 2136 94 2141 97
rect 2143 105 2150 107
rect 2143 103 2146 105
rect 2148 103 2150 105
rect 2143 101 2150 103
rect 2155 101 2160 108
rect 2176 105 2182 108
rect 2184 112 2191 114
rect 2184 110 2187 112
rect 2189 110 2191 112
rect 2184 108 2191 110
rect 2245 108 2250 109
rect 2184 105 2189 108
rect 2199 106 2206 108
rect 2176 101 2180 105
rect 2143 94 2148 101
rect 2155 99 2161 101
rect 2155 97 2157 99
rect 2159 97 2161 99
rect 2155 95 2161 97
rect 2174 99 2180 101
rect 2199 104 2201 106
rect 2203 104 2206 106
rect 2199 102 2206 104
rect 2208 106 2216 108
rect 2208 104 2211 106
rect 2213 104 2216 106
rect 2208 102 2216 104
rect 2174 97 2176 99
rect 2178 97 2180 99
rect 2174 95 2180 97
rect 2210 100 2216 102
rect 2218 100 2223 108
rect 2225 104 2233 108
rect 2225 102 2228 104
rect 2230 102 2233 104
rect 2225 100 2233 102
rect 2235 100 2240 108
rect 2242 104 2250 108
rect 2242 102 2245 104
rect 2247 102 2250 104
rect 2242 100 2250 102
rect 2252 107 2259 109
rect 2313 108 2318 109
rect 2252 105 2255 107
rect 2257 105 2259 107
rect 2252 103 2259 105
rect 2267 106 2274 108
rect 2267 104 2269 106
rect 2271 104 2274 106
rect 2252 100 2257 103
rect 2267 102 2274 104
rect 2276 106 2284 108
rect 2276 104 2279 106
rect 2281 104 2284 106
rect 2276 102 2284 104
rect 2278 100 2284 102
rect 2286 100 2291 108
rect 2293 104 2301 108
rect 2293 102 2296 104
rect 2298 102 2301 104
rect 2293 100 2301 102
rect 2303 100 2308 108
rect 2310 104 2318 108
rect 2310 102 2313 104
rect 2315 102 2318 104
rect 2310 100 2318 102
rect 2320 107 2327 109
rect 2320 105 2323 107
rect 2325 105 2327 107
rect 2320 103 2327 105
rect 2320 100 2325 103
rect 26 83 33 85
rect 26 81 29 83
rect 31 81 33 83
rect 26 75 33 81
rect 66 83 73 85
rect 66 81 69 83
rect 71 81 73 83
rect 8 73 15 75
rect 8 71 10 73
rect 12 71 15 73
rect 8 69 15 71
rect 10 64 15 69
rect 17 64 22 75
rect 24 73 33 75
rect 66 75 73 81
rect 48 73 55 75
rect 24 64 35 73
rect 37 71 44 73
rect 37 69 40 71
rect 42 69 44 71
rect 48 71 50 73
rect 52 71 55 73
rect 48 69 55 71
rect 37 67 44 69
rect 37 64 42 67
rect 50 64 55 69
rect 57 64 62 75
rect 64 73 73 75
rect 90 75 95 82
rect 88 73 95 75
rect 64 64 75 73
rect 77 71 84 73
rect 77 69 80 71
rect 82 69 84 71
rect 88 71 90 73
rect 92 71 95 73
rect 88 69 95 71
rect 97 79 102 82
rect 97 77 105 79
rect 97 75 100 77
rect 102 75 105 77
rect 97 69 105 75
rect 107 76 112 79
rect 107 74 115 76
rect 107 72 110 74
rect 112 72 115 74
rect 107 69 115 72
rect 77 67 84 69
rect 77 64 82 67
rect 110 62 115 69
rect 117 66 125 76
rect 117 64 120 66
rect 122 64 125 66
rect 117 62 125 64
rect 127 73 134 76
rect 140 75 145 82
rect 127 71 130 73
rect 132 71 134 73
rect 127 66 134 71
rect 138 73 145 75
rect 138 71 140 73
rect 142 71 145 73
rect 138 69 145 71
rect 127 64 130 66
rect 132 64 134 66
rect 127 62 134 64
rect 140 62 145 69
rect 147 62 152 82
rect 154 80 163 82
rect 154 78 157 80
rect 159 78 163 80
rect 154 68 163 78
rect 165 75 170 82
rect 180 75 185 82
rect 165 73 172 75
rect 165 71 168 73
rect 170 71 172 73
rect 165 68 172 71
rect 178 73 185 75
rect 178 71 180 73
rect 182 71 185 73
rect 178 68 185 71
rect 187 80 196 82
rect 187 78 191 80
rect 193 78 196 80
rect 187 68 196 78
rect 154 62 161 68
rect 189 62 196 68
rect 198 62 203 82
rect 205 75 210 82
rect 248 79 253 82
rect 238 76 243 79
rect 205 73 212 75
rect 205 71 208 73
rect 210 71 212 73
rect 205 69 212 71
rect 216 73 223 76
rect 216 71 218 73
rect 220 71 223 73
rect 205 62 210 69
rect 216 66 223 71
rect 216 64 218 66
rect 220 64 223 66
rect 216 62 223 64
rect 225 66 233 76
rect 225 64 228 66
rect 230 64 233 66
rect 225 62 233 64
rect 235 74 243 76
rect 235 72 238 74
rect 240 72 243 74
rect 235 69 243 72
rect 245 77 253 79
rect 245 75 248 77
rect 250 75 253 77
rect 245 69 253 75
rect 255 75 260 82
rect 267 79 273 81
rect 267 77 269 79
rect 271 77 273 79
rect 267 75 273 77
rect 286 79 292 81
rect 333 83 340 85
rect 333 81 336 83
rect 338 81 340 83
rect 286 77 288 79
rect 290 77 292 79
rect 286 75 292 77
rect 255 73 262 75
rect 255 71 258 73
rect 260 71 262 73
rect 255 69 262 71
rect 235 62 240 69
rect 267 68 272 75
rect 288 71 292 75
rect 333 75 340 81
rect 315 73 322 75
rect 315 71 317 73
rect 319 71 322 73
rect 288 68 294 71
rect 267 62 274 68
rect 276 66 284 68
rect 276 64 279 66
rect 281 64 284 66
rect 276 62 284 64
rect 286 62 294 68
rect 296 68 301 71
rect 315 69 322 71
rect 296 66 303 68
rect 296 64 299 66
rect 301 64 303 66
rect 317 64 322 69
rect 324 64 329 75
rect 331 73 340 75
rect 357 75 362 82
rect 355 73 362 75
rect 331 64 342 73
rect 344 71 351 73
rect 344 69 347 71
rect 349 69 351 71
rect 355 71 357 73
rect 359 71 362 73
rect 355 69 362 71
rect 364 79 369 82
rect 364 77 372 79
rect 364 75 367 77
rect 369 75 372 77
rect 364 69 372 75
rect 374 76 379 79
rect 374 74 382 76
rect 374 72 377 74
rect 379 72 382 74
rect 374 69 382 72
rect 344 67 351 69
rect 344 64 349 67
rect 296 62 303 64
rect 377 62 382 69
rect 384 66 392 76
rect 384 64 387 66
rect 389 64 392 66
rect 384 62 392 64
rect 394 73 401 76
rect 407 75 412 82
rect 394 71 397 73
rect 399 71 401 73
rect 394 66 401 71
rect 405 73 412 75
rect 405 71 407 73
rect 409 71 412 73
rect 405 69 412 71
rect 394 64 397 66
rect 399 64 401 66
rect 394 62 401 64
rect 407 62 412 69
rect 414 62 419 82
rect 421 80 430 82
rect 421 78 424 80
rect 426 78 430 80
rect 421 68 430 78
rect 432 75 437 82
rect 447 75 452 82
rect 432 73 439 75
rect 432 71 435 73
rect 437 71 439 73
rect 432 68 439 71
rect 445 73 452 75
rect 445 71 447 73
rect 449 71 452 73
rect 445 68 452 71
rect 454 80 463 82
rect 454 78 458 80
rect 460 78 463 80
rect 454 68 463 78
rect 421 62 428 68
rect 456 62 463 68
rect 465 62 470 82
rect 472 75 477 82
rect 515 79 520 82
rect 505 76 510 79
rect 472 73 479 75
rect 472 71 475 73
rect 477 71 479 73
rect 472 69 479 71
rect 483 73 490 76
rect 483 71 485 73
rect 487 71 490 73
rect 472 62 477 69
rect 483 66 490 71
rect 483 64 485 66
rect 487 64 490 66
rect 483 62 490 64
rect 492 66 500 76
rect 492 64 495 66
rect 497 64 500 66
rect 492 62 500 64
rect 502 74 510 76
rect 502 72 505 74
rect 507 72 510 74
rect 502 69 510 72
rect 512 77 520 79
rect 512 75 515 77
rect 517 75 520 77
rect 512 69 520 75
rect 522 75 527 82
rect 534 79 540 81
rect 534 77 536 79
rect 538 77 540 79
rect 534 75 540 77
rect 553 79 559 81
rect 600 83 607 85
rect 600 81 603 83
rect 605 81 607 83
rect 553 77 555 79
rect 557 77 559 79
rect 553 75 559 77
rect 522 73 529 75
rect 522 71 525 73
rect 527 71 529 73
rect 522 69 529 71
rect 502 62 507 69
rect 534 68 539 75
rect 555 71 559 75
rect 600 75 607 81
rect 582 73 589 75
rect 582 71 584 73
rect 586 71 589 73
rect 555 68 561 71
rect 534 62 541 68
rect 543 66 551 68
rect 543 64 546 66
rect 548 64 551 66
rect 543 62 551 64
rect 553 62 561 68
rect 563 68 568 71
rect 582 69 589 71
rect 563 66 570 68
rect 563 64 566 66
rect 568 64 570 66
rect 584 64 589 69
rect 591 64 596 75
rect 598 73 607 75
rect 624 75 629 82
rect 622 73 629 75
rect 598 64 609 73
rect 611 71 618 73
rect 611 69 614 71
rect 616 69 618 71
rect 622 71 624 73
rect 626 71 629 73
rect 622 69 629 71
rect 631 79 636 82
rect 631 77 639 79
rect 631 75 634 77
rect 636 75 639 77
rect 631 69 639 75
rect 641 76 646 79
rect 641 74 649 76
rect 641 72 644 74
rect 646 72 649 74
rect 641 69 649 72
rect 611 67 618 69
rect 611 64 616 67
rect 563 62 570 64
rect 644 62 649 69
rect 651 66 659 76
rect 651 64 654 66
rect 656 64 659 66
rect 651 62 659 64
rect 661 73 668 76
rect 674 75 679 82
rect 661 71 664 73
rect 666 71 668 73
rect 661 66 668 71
rect 672 73 679 75
rect 672 71 674 73
rect 676 71 679 73
rect 672 69 679 71
rect 661 64 664 66
rect 666 64 668 66
rect 661 62 668 64
rect 674 62 679 69
rect 681 62 686 82
rect 688 80 697 82
rect 688 78 691 80
rect 693 78 697 80
rect 688 68 697 78
rect 699 75 704 82
rect 714 75 719 82
rect 699 73 706 75
rect 699 71 702 73
rect 704 71 706 73
rect 699 68 706 71
rect 712 73 719 75
rect 712 71 714 73
rect 716 71 719 73
rect 712 68 719 71
rect 721 80 730 82
rect 721 78 725 80
rect 727 78 730 80
rect 721 68 730 78
rect 688 62 695 68
rect 723 62 730 68
rect 732 62 737 82
rect 739 75 744 82
rect 782 79 787 82
rect 772 76 777 79
rect 739 73 746 75
rect 739 71 742 73
rect 744 71 746 73
rect 739 69 746 71
rect 750 73 757 76
rect 750 71 752 73
rect 754 71 757 73
rect 739 62 744 69
rect 750 66 757 71
rect 750 64 752 66
rect 754 64 757 66
rect 750 62 757 64
rect 759 66 767 76
rect 759 64 762 66
rect 764 64 767 66
rect 759 62 767 64
rect 769 74 777 76
rect 769 72 772 74
rect 774 72 777 74
rect 769 69 777 72
rect 779 77 787 79
rect 779 75 782 77
rect 784 75 787 77
rect 779 69 787 75
rect 789 75 794 82
rect 801 79 807 81
rect 801 77 803 79
rect 805 77 807 79
rect 801 75 807 77
rect 820 79 826 81
rect 867 83 874 85
rect 867 81 870 83
rect 872 81 874 83
rect 820 77 822 79
rect 824 77 826 79
rect 820 75 826 77
rect 789 73 796 75
rect 789 71 792 73
rect 794 71 796 73
rect 789 69 796 71
rect 769 62 774 69
rect 801 68 806 75
rect 822 71 826 75
rect 867 75 874 81
rect 849 73 856 75
rect 849 71 851 73
rect 853 71 856 73
rect 822 68 828 71
rect 801 62 808 68
rect 810 66 818 68
rect 810 64 813 66
rect 815 64 818 66
rect 810 62 818 64
rect 820 62 828 68
rect 830 68 835 71
rect 849 69 856 71
rect 830 66 837 68
rect 830 64 833 66
rect 835 64 837 66
rect 851 64 856 69
rect 858 64 863 75
rect 865 73 874 75
rect 891 75 896 82
rect 889 73 896 75
rect 865 64 876 73
rect 878 71 885 73
rect 878 69 881 71
rect 883 69 885 71
rect 889 71 891 73
rect 893 71 896 73
rect 889 69 896 71
rect 898 79 903 82
rect 898 77 906 79
rect 898 75 901 77
rect 903 75 906 77
rect 898 69 906 75
rect 908 76 913 79
rect 908 74 916 76
rect 908 72 911 74
rect 913 72 916 74
rect 908 69 916 72
rect 878 67 885 69
rect 878 64 883 67
rect 830 62 837 64
rect 911 62 916 69
rect 918 66 926 76
rect 918 64 921 66
rect 923 64 926 66
rect 918 62 926 64
rect 928 73 935 76
rect 941 75 946 82
rect 928 71 931 73
rect 933 71 935 73
rect 928 66 935 71
rect 939 73 946 75
rect 939 71 941 73
rect 943 71 946 73
rect 939 69 946 71
rect 928 64 931 66
rect 933 64 935 66
rect 928 62 935 64
rect 941 62 946 69
rect 948 62 953 82
rect 955 80 964 82
rect 955 78 958 80
rect 960 78 964 80
rect 955 68 964 78
rect 966 75 971 82
rect 981 75 986 82
rect 966 73 973 75
rect 966 71 969 73
rect 971 71 973 73
rect 966 68 973 71
rect 979 73 986 75
rect 979 71 981 73
rect 983 71 986 73
rect 979 68 986 71
rect 988 80 997 82
rect 988 78 992 80
rect 994 78 997 80
rect 988 68 997 78
rect 955 62 962 68
rect 990 62 997 68
rect 999 62 1004 82
rect 1006 75 1011 82
rect 1049 79 1054 82
rect 1039 76 1044 79
rect 1006 73 1013 75
rect 1006 71 1009 73
rect 1011 71 1013 73
rect 1006 69 1013 71
rect 1017 73 1024 76
rect 1017 71 1019 73
rect 1021 71 1024 73
rect 1006 62 1011 69
rect 1017 66 1024 71
rect 1017 64 1019 66
rect 1021 64 1024 66
rect 1017 62 1024 64
rect 1026 66 1034 76
rect 1026 64 1029 66
rect 1031 64 1034 66
rect 1026 62 1034 64
rect 1036 74 1044 76
rect 1036 72 1039 74
rect 1041 72 1044 74
rect 1036 69 1044 72
rect 1046 77 1054 79
rect 1046 75 1049 77
rect 1051 75 1054 77
rect 1046 69 1054 75
rect 1056 75 1061 82
rect 1068 79 1074 81
rect 1068 77 1070 79
rect 1072 77 1074 79
rect 1068 75 1074 77
rect 1087 79 1093 81
rect 1134 83 1141 85
rect 1134 81 1137 83
rect 1139 81 1141 83
rect 1087 77 1089 79
rect 1091 77 1093 79
rect 1087 75 1093 77
rect 1056 73 1063 75
rect 1056 71 1059 73
rect 1061 71 1063 73
rect 1056 69 1063 71
rect 1036 62 1041 69
rect 1068 68 1073 75
rect 1089 71 1093 75
rect 1134 75 1141 81
rect 1116 73 1123 75
rect 1116 71 1118 73
rect 1120 71 1123 73
rect 1089 68 1095 71
rect 1068 62 1075 68
rect 1077 66 1085 68
rect 1077 64 1080 66
rect 1082 64 1085 66
rect 1077 62 1085 64
rect 1087 62 1095 68
rect 1097 68 1102 71
rect 1116 69 1123 71
rect 1097 66 1104 68
rect 1097 64 1100 66
rect 1102 64 1104 66
rect 1118 64 1123 69
rect 1125 64 1130 75
rect 1132 73 1141 75
rect 1158 75 1163 82
rect 1156 73 1163 75
rect 1132 64 1143 73
rect 1145 71 1152 73
rect 1145 69 1148 71
rect 1150 69 1152 71
rect 1156 71 1158 73
rect 1160 71 1163 73
rect 1156 69 1163 71
rect 1165 79 1170 82
rect 1165 77 1173 79
rect 1165 75 1168 77
rect 1170 75 1173 77
rect 1165 69 1173 75
rect 1175 76 1180 79
rect 1175 74 1183 76
rect 1175 72 1178 74
rect 1180 72 1183 74
rect 1175 69 1183 72
rect 1145 67 1152 69
rect 1145 64 1150 67
rect 1097 62 1104 64
rect 1178 62 1183 69
rect 1185 66 1193 76
rect 1185 64 1188 66
rect 1190 64 1193 66
rect 1185 62 1193 64
rect 1195 73 1202 76
rect 1208 75 1213 82
rect 1195 71 1198 73
rect 1200 71 1202 73
rect 1195 66 1202 71
rect 1206 73 1213 75
rect 1206 71 1208 73
rect 1210 71 1213 73
rect 1206 69 1213 71
rect 1195 64 1198 66
rect 1200 64 1202 66
rect 1195 62 1202 64
rect 1208 62 1213 69
rect 1215 62 1220 82
rect 1222 80 1231 82
rect 1222 78 1225 80
rect 1227 78 1231 80
rect 1222 68 1231 78
rect 1233 75 1238 82
rect 1248 75 1253 82
rect 1233 73 1240 75
rect 1233 71 1236 73
rect 1238 71 1240 73
rect 1233 68 1240 71
rect 1246 73 1253 75
rect 1246 71 1248 73
rect 1250 71 1253 73
rect 1246 68 1253 71
rect 1255 80 1264 82
rect 1255 78 1259 80
rect 1261 78 1264 80
rect 1255 68 1264 78
rect 1222 62 1229 68
rect 1257 62 1264 68
rect 1266 62 1271 82
rect 1273 75 1278 82
rect 1316 79 1321 82
rect 1306 76 1311 79
rect 1273 73 1280 75
rect 1273 71 1276 73
rect 1278 71 1280 73
rect 1273 69 1280 71
rect 1284 73 1291 76
rect 1284 71 1286 73
rect 1288 71 1291 73
rect 1273 62 1278 69
rect 1284 66 1291 71
rect 1284 64 1286 66
rect 1288 64 1291 66
rect 1284 62 1291 64
rect 1293 66 1301 76
rect 1293 64 1296 66
rect 1298 64 1301 66
rect 1293 62 1301 64
rect 1303 74 1311 76
rect 1303 72 1306 74
rect 1308 72 1311 74
rect 1303 69 1311 72
rect 1313 77 1321 79
rect 1313 75 1316 77
rect 1318 75 1321 77
rect 1313 69 1321 75
rect 1323 75 1328 82
rect 1335 79 1341 81
rect 1335 77 1337 79
rect 1339 77 1341 79
rect 1335 75 1341 77
rect 1354 79 1360 81
rect 1401 83 1408 85
rect 1401 81 1404 83
rect 1406 81 1408 83
rect 1354 77 1356 79
rect 1358 77 1360 79
rect 1354 75 1360 77
rect 1323 73 1330 75
rect 1323 71 1326 73
rect 1328 71 1330 73
rect 1323 69 1330 71
rect 1303 62 1308 69
rect 1335 68 1340 75
rect 1356 71 1360 75
rect 1401 75 1408 81
rect 1383 73 1390 75
rect 1383 71 1385 73
rect 1387 71 1390 73
rect 1356 68 1362 71
rect 1335 62 1342 68
rect 1344 66 1352 68
rect 1344 64 1347 66
rect 1349 64 1352 66
rect 1344 62 1352 64
rect 1354 62 1362 68
rect 1364 68 1369 71
rect 1383 69 1390 71
rect 1364 66 1371 68
rect 1364 64 1367 66
rect 1369 64 1371 66
rect 1385 64 1390 69
rect 1392 64 1397 75
rect 1399 73 1408 75
rect 1425 75 1430 82
rect 1423 73 1430 75
rect 1399 64 1410 73
rect 1412 71 1419 73
rect 1412 69 1415 71
rect 1417 69 1419 71
rect 1423 71 1425 73
rect 1427 71 1430 73
rect 1423 69 1430 71
rect 1432 79 1437 82
rect 1432 77 1440 79
rect 1432 75 1435 77
rect 1437 75 1440 77
rect 1432 69 1440 75
rect 1442 76 1447 79
rect 1442 74 1450 76
rect 1442 72 1445 74
rect 1447 72 1450 74
rect 1442 69 1450 72
rect 1412 67 1419 69
rect 1412 64 1417 67
rect 1364 62 1371 64
rect 1445 62 1450 69
rect 1452 66 1460 76
rect 1452 64 1455 66
rect 1457 64 1460 66
rect 1452 62 1460 64
rect 1462 73 1469 76
rect 1475 75 1480 82
rect 1462 71 1465 73
rect 1467 71 1469 73
rect 1462 66 1469 71
rect 1473 73 1480 75
rect 1473 71 1475 73
rect 1477 71 1480 73
rect 1473 69 1480 71
rect 1462 64 1465 66
rect 1467 64 1469 66
rect 1462 62 1469 64
rect 1475 62 1480 69
rect 1482 62 1487 82
rect 1489 80 1498 82
rect 1489 78 1492 80
rect 1494 78 1498 80
rect 1489 68 1498 78
rect 1500 75 1505 82
rect 1515 75 1520 82
rect 1500 73 1507 75
rect 1500 71 1503 73
rect 1505 71 1507 73
rect 1500 68 1507 71
rect 1513 73 1520 75
rect 1513 71 1515 73
rect 1517 71 1520 73
rect 1513 68 1520 71
rect 1522 80 1531 82
rect 1522 78 1526 80
rect 1528 78 1531 80
rect 1522 68 1531 78
rect 1489 62 1496 68
rect 1524 62 1531 68
rect 1533 62 1538 82
rect 1540 75 1545 82
rect 1583 79 1588 82
rect 1573 76 1578 79
rect 1540 73 1547 75
rect 1540 71 1543 73
rect 1545 71 1547 73
rect 1540 69 1547 71
rect 1551 73 1558 76
rect 1551 71 1553 73
rect 1555 71 1558 73
rect 1540 62 1545 69
rect 1551 66 1558 71
rect 1551 64 1553 66
rect 1555 64 1558 66
rect 1551 62 1558 64
rect 1560 66 1568 76
rect 1560 64 1563 66
rect 1565 64 1568 66
rect 1560 62 1568 64
rect 1570 74 1578 76
rect 1570 72 1573 74
rect 1575 72 1578 74
rect 1570 69 1578 72
rect 1580 77 1588 79
rect 1580 75 1583 77
rect 1585 75 1588 77
rect 1580 69 1588 75
rect 1590 75 1595 82
rect 1602 79 1608 81
rect 1602 77 1604 79
rect 1606 77 1608 79
rect 1602 75 1608 77
rect 1621 79 1627 81
rect 1668 83 1675 85
rect 1668 81 1671 83
rect 1673 81 1675 83
rect 1621 77 1623 79
rect 1625 77 1627 79
rect 1621 75 1627 77
rect 1590 73 1597 75
rect 1590 71 1593 73
rect 1595 71 1597 73
rect 1590 69 1597 71
rect 1570 62 1575 69
rect 1602 68 1607 75
rect 1623 71 1627 75
rect 1668 75 1675 81
rect 1650 73 1657 75
rect 1650 71 1652 73
rect 1654 71 1657 73
rect 1623 68 1629 71
rect 1602 62 1609 68
rect 1611 66 1619 68
rect 1611 64 1614 66
rect 1616 64 1619 66
rect 1611 62 1619 64
rect 1621 62 1629 68
rect 1631 68 1636 71
rect 1650 69 1657 71
rect 1631 66 1638 68
rect 1631 64 1634 66
rect 1636 64 1638 66
rect 1652 64 1657 69
rect 1659 64 1664 75
rect 1666 73 1675 75
rect 1692 75 1697 82
rect 1690 73 1697 75
rect 1666 64 1677 73
rect 1679 71 1686 73
rect 1679 69 1682 71
rect 1684 69 1686 71
rect 1690 71 1692 73
rect 1694 71 1697 73
rect 1690 69 1697 71
rect 1699 79 1704 82
rect 1699 77 1707 79
rect 1699 75 1702 77
rect 1704 75 1707 77
rect 1699 69 1707 75
rect 1709 76 1714 79
rect 1709 74 1717 76
rect 1709 72 1712 74
rect 1714 72 1717 74
rect 1709 69 1717 72
rect 1679 67 1686 69
rect 1679 64 1684 67
rect 1631 62 1638 64
rect 1712 62 1717 69
rect 1719 66 1727 76
rect 1719 64 1722 66
rect 1724 64 1727 66
rect 1719 62 1727 64
rect 1729 73 1736 76
rect 1742 75 1747 82
rect 1729 71 1732 73
rect 1734 71 1736 73
rect 1729 66 1736 71
rect 1740 73 1747 75
rect 1740 71 1742 73
rect 1744 71 1747 73
rect 1740 69 1747 71
rect 1729 64 1732 66
rect 1734 64 1736 66
rect 1729 62 1736 64
rect 1742 62 1747 69
rect 1749 62 1754 82
rect 1756 80 1765 82
rect 1756 78 1759 80
rect 1761 78 1765 80
rect 1756 68 1765 78
rect 1767 75 1772 82
rect 1782 75 1787 82
rect 1767 73 1774 75
rect 1767 71 1770 73
rect 1772 71 1774 73
rect 1767 68 1774 71
rect 1780 73 1787 75
rect 1780 71 1782 73
rect 1784 71 1787 73
rect 1780 68 1787 71
rect 1789 80 1798 82
rect 1789 78 1793 80
rect 1795 78 1798 80
rect 1789 68 1798 78
rect 1756 62 1763 68
rect 1791 62 1798 68
rect 1800 62 1805 82
rect 1807 75 1812 82
rect 1850 79 1855 82
rect 1840 76 1845 79
rect 1807 73 1814 75
rect 1807 71 1810 73
rect 1812 71 1814 73
rect 1807 69 1814 71
rect 1818 73 1825 76
rect 1818 71 1820 73
rect 1822 71 1825 73
rect 1807 62 1812 69
rect 1818 66 1825 71
rect 1818 64 1820 66
rect 1822 64 1825 66
rect 1818 62 1825 64
rect 1827 66 1835 76
rect 1827 64 1830 66
rect 1832 64 1835 66
rect 1827 62 1835 64
rect 1837 74 1845 76
rect 1837 72 1840 74
rect 1842 72 1845 74
rect 1837 69 1845 72
rect 1847 77 1855 79
rect 1847 75 1850 77
rect 1852 75 1855 77
rect 1847 69 1855 75
rect 1857 75 1862 82
rect 1869 79 1875 81
rect 1869 77 1871 79
rect 1873 77 1875 79
rect 1869 75 1875 77
rect 1888 79 1894 81
rect 1888 77 1890 79
rect 1892 77 1894 79
rect 1888 75 1894 77
rect 1966 83 1972 85
rect 1966 81 1968 83
rect 1970 81 1972 83
rect 1966 79 1972 81
rect 1950 76 1955 79
rect 1857 73 1864 75
rect 1857 71 1860 73
rect 1862 71 1864 73
rect 1857 69 1864 71
rect 1837 62 1842 69
rect 1869 68 1874 75
rect 1890 71 1894 75
rect 1926 74 1935 76
rect 1926 72 1928 74
rect 1930 72 1935 74
rect 1926 71 1935 72
rect 1890 68 1896 71
rect 1869 62 1876 68
rect 1878 66 1886 68
rect 1878 64 1881 66
rect 1883 64 1886 66
rect 1878 62 1886 64
rect 1888 62 1896 68
rect 1898 68 1903 71
rect 1914 68 1919 71
rect 1898 66 1905 68
rect 1898 64 1901 66
rect 1903 64 1905 66
rect 1898 62 1905 64
rect 1912 66 1919 68
rect 1912 64 1914 66
rect 1916 64 1919 66
rect 1912 62 1919 64
rect 1921 67 1935 71
rect 1937 71 1945 76
rect 1937 69 1940 71
rect 1942 69 1945 71
rect 1937 67 1945 69
rect 1947 73 1955 76
rect 1947 71 1950 73
rect 1952 71 1955 73
rect 1947 67 1955 71
rect 1957 67 1962 79
rect 1964 67 1972 79
rect 1978 75 1983 82
rect 1976 73 1983 75
rect 1976 71 1978 73
rect 1980 71 1983 73
rect 1976 69 1983 71
rect 1985 79 1990 82
rect 1985 77 1993 79
rect 1985 75 1988 77
rect 1990 75 1993 77
rect 1985 69 1993 75
rect 1995 76 2000 79
rect 1995 74 2003 76
rect 1995 72 1998 74
rect 2000 72 2003 74
rect 1995 69 2003 72
rect 1921 62 1926 67
rect 1998 62 2003 69
rect 2005 66 2013 76
rect 2005 64 2008 66
rect 2010 64 2013 66
rect 2005 62 2013 64
rect 2015 73 2022 76
rect 2028 75 2033 82
rect 2015 71 2018 73
rect 2020 71 2022 73
rect 2015 66 2022 71
rect 2026 73 2033 75
rect 2026 71 2028 73
rect 2030 71 2033 73
rect 2026 69 2033 71
rect 2015 64 2018 66
rect 2020 64 2022 66
rect 2015 62 2022 64
rect 2028 62 2033 69
rect 2035 62 2040 82
rect 2042 80 2051 82
rect 2042 78 2045 80
rect 2047 78 2051 80
rect 2042 68 2051 78
rect 2053 75 2058 82
rect 2068 75 2073 82
rect 2053 73 2060 75
rect 2053 71 2056 73
rect 2058 71 2060 73
rect 2053 68 2060 71
rect 2066 73 2073 75
rect 2066 71 2068 73
rect 2070 71 2073 73
rect 2066 68 2073 71
rect 2075 80 2084 82
rect 2075 78 2079 80
rect 2081 78 2084 80
rect 2075 68 2084 78
rect 2042 62 2049 68
rect 2077 62 2084 68
rect 2086 62 2091 82
rect 2093 75 2098 82
rect 2136 79 2141 82
rect 2126 76 2131 79
rect 2093 73 2100 75
rect 2093 71 2096 73
rect 2098 71 2100 73
rect 2093 69 2100 71
rect 2104 73 2111 76
rect 2104 71 2106 73
rect 2108 71 2111 73
rect 2093 62 2098 69
rect 2104 66 2111 71
rect 2104 64 2106 66
rect 2108 64 2111 66
rect 2104 62 2111 64
rect 2113 66 2121 76
rect 2113 64 2116 66
rect 2118 64 2121 66
rect 2113 62 2121 64
rect 2123 74 2131 76
rect 2123 72 2126 74
rect 2128 72 2131 74
rect 2123 69 2131 72
rect 2133 77 2141 79
rect 2133 75 2136 77
rect 2138 75 2141 77
rect 2133 69 2141 75
rect 2143 75 2148 82
rect 2155 79 2161 81
rect 2155 77 2157 79
rect 2159 77 2161 79
rect 2155 75 2161 77
rect 2174 79 2180 81
rect 2174 77 2176 79
rect 2178 77 2180 79
rect 2174 75 2180 77
rect 2143 73 2150 75
rect 2143 71 2146 73
rect 2148 71 2150 73
rect 2143 69 2150 71
rect 2123 62 2128 69
rect 2155 68 2160 75
rect 2176 71 2180 75
rect 2210 74 2216 76
rect 2199 72 2206 74
rect 2176 68 2182 71
rect 2155 62 2162 68
rect 2164 66 2172 68
rect 2164 64 2167 66
rect 2169 64 2172 66
rect 2164 62 2172 64
rect 2174 62 2182 68
rect 2184 68 2189 71
rect 2199 70 2201 72
rect 2203 70 2206 72
rect 2199 68 2206 70
rect 2208 72 2216 74
rect 2208 70 2211 72
rect 2213 70 2216 72
rect 2208 68 2216 70
rect 2218 68 2223 76
rect 2225 74 2233 76
rect 2225 72 2228 74
rect 2230 72 2233 74
rect 2225 68 2233 72
rect 2235 68 2240 76
rect 2242 74 2250 76
rect 2242 72 2245 74
rect 2247 72 2250 74
rect 2242 68 2250 72
rect 2184 66 2191 68
rect 2184 64 2187 66
rect 2189 64 2191 66
rect 2184 62 2191 64
rect 2245 67 2250 68
rect 2252 73 2257 76
rect 2278 74 2284 76
rect 2252 71 2259 73
rect 2252 69 2255 71
rect 2257 69 2259 71
rect 2252 67 2259 69
rect 2267 72 2274 74
rect 2267 70 2269 72
rect 2271 70 2274 72
rect 2267 68 2274 70
rect 2276 72 2284 74
rect 2276 70 2279 72
rect 2281 70 2284 72
rect 2276 68 2284 70
rect 2286 68 2291 76
rect 2293 74 2301 76
rect 2293 72 2296 74
rect 2298 72 2301 74
rect 2293 68 2301 72
rect 2303 68 2308 76
rect 2310 74 2318 76
rect 2310 72 2313 74
rect 2315 72 2318 74
rect 2310 68 2318 72
rect 2313 67 2318 68
rect 2320 73 2325 76
rect 2320 71 2327 73
rect 2320 69 2323 71
rect 2325 69 2327 71
rect 2320 67 2327 69
rect 10 -37 15 -32
rect 8 -39 15 -37
rect 8 -41 10 -39
rect 12 -41 15 -39
rect 8 -43 15 -41
rect 17 -43 22 -32
rect 24 -41 35 -32
rect 37 -35 42 -32
rect 37 -37 44 -35
rect 50 -37 55 -32
rect 37 -39 40 -37
rect 42 -39 44 -37
rect 37 -41 44 -39
rect 48 -39 55 -37
rect 48 -41 50 -39
rect 52 -41 55 -39
rect 24 -43 33 -41
rect 26 -49 33 -43
rect 48 -43 55 -41
rect 57 -43 62 -32
rect 64 -41 75 -32
rect 77 -35 82 -32
rect 77 -37 84 -35
rect 110 -37 115 -30
rect 77 -39 80 -37
rect 82 -39 84 -37
rect 77 -41 84 -39
rect 88 -39 95 -37
rect 88 -41 90 -39
rect 92 -41 95 -39
rect 64 -43 73 -41
rect 26 -51 29 -49
rect 31 -51 33 -49
rect 26 -53 33 -51
rect 66 -49 73 -43
rect 88 -43 95 -41
rect 66 -51 69 -49
rect 71 -51 73 -49
rect 66 -53 73 -51
rect 90 -50 95 -43
rect 97 -43 105 -37
rect 97 -45 100 -43
rect 102 -45 105 -43
rect 97 -47 105 -45
rect 107 -40 115 -37
rect 107 -42 110 -40
rect 112 -42 115 -40
rect 107 -44 115 -42
rect 117 -32 125 -30
rect 117 -34 120 -32
rect 122 -34 125 -32
rect 117 -44 125 -34
rect 127 -32 134 -30
rect 127 -34 130 -32
rect 132 -34 134 -32
rect 127 -39 134 -34
rect 140 -37 145 -30
rect 127 -41 130 -39
rect 132 -41 134 -39
rect 127 -44 134 -41
rect 138 -39 145 -37
rect 138 -41 140 -39
rect 142 -41 145 -39
rect 138 -43 145 -41
rect 107 -47 112 -44
rect 97 -50 102 -47
rect 140 -50 145 -43
rect 147 -50 152 -30
rect 154 -36 161 -30
rect 189 -36 196 -30
rect 154 -46 163 -36
rect 154 -48 157 -46
rect 159 -48 163 -46
rect 154 -50 163 -48
rect 165 -39 172 -36
rect 165 -41 168 -39
rect 170 -41 172 -39
rect 165 -43 172 -41
rect 178 -39 185 -36
rect 178 -41 180 -39
rect 182 -41 185 -39
rect 178 -43 185 -41
rect 165 -50 170 -43
rect 180 -50 185 -43
rect 187 -46 196 -36
rect 187 -48 191 -46
rect 193 -48 196 -46
rect 187 -50 196 -48
rect 198 -50 203 -30
rect 205 -37 210 -30
rect 216 -32 223 -30
rect 216 -34 218 -32
rect 220 -34 223 -32
rect 205 -39 212 -37
rect 205 -41 208 -39
rect 210 -41 212 -39
rect 205 -43 212 -41
rect 216 -39 223 -34
rect 216 -41 218 -39
rect 220 -41 223 -39
rect 205 -50 210 -43
rect 216 -44 223 -41
rect 225 -32 233 -30
rect 225 -34 228 -32
rect 230 -34 233 -32
rect 225 -44 233 -34
rect 235 -37 240 -30
rect 267 -36 274 -30
rect 276 -32 284 -30
rect 276 -34 279 -32
rect 281 -34 284 -32
rect 276 -36 284 -34
rect 286 -36 294 -30
rect 235 -40 243 -37
rect 235 -42 238 -40
rect 240 -42 243 -40
rect 235 -44 243 -42
rect 238 -47 243 -44
rect 245 -43 253 -37
rect 245 -45 248 -43
rect 250 -45 253 -43
rect 245 -47 253 -45
rect 248 -50 253 -47
rect 255 -39 262 -37
rect 255 -41 258 -39
rect 260 -41 262 -39
rect 255 -43 262 -41
rect 267 -43 272 -36
rect 288 -39 294 -36
rect 296 -32 303 -30
rect 296 -34 299 -32
rect 301 -34 303 -32
rect 296 -36 303 -34
rect 296 -39 301 -36
rect 317 -37 322 -32
rect 315 -39 322 -37
rect 288 -43 292 -39
rect 255 -50 260 -43
rect 267 -45 273 -43
rect 267 -47 269 -45
rect 271 -47 273 -45
rect 267 -49 273 -47
rect 286 -45 292 -43
rect 315 -41 317 -39
rect 319 -41 322 -39
rect 315 -43 322 -41
rect 324 -43 329 -32
rect 331 -41 342 -32
rect 344 -35 349 -32
rect 344 -37 351 -35
rect 377 -37 382 -30
rect 344 -39 347 -37
rect 349 -39 351 -37
rect 344 -41 351 -39
rect 355 -39 362 -37
rect 355 -41 357 -39
rect 359 -41 362 -39
rect 331 -43 340 -41
rect 286 -47 288 -45
rect 290 -47 292 -45
rect 286 -49 292 -47
rect 333 -49 340 -43
rect 355 -43 362 -41
rect 333 -51 336 -49
rect 338 -51 340 -49
rect 333 -53 340 -51
rect 357 -50 362 -43
rect 364 -43 372 -37
rect 364 -45 367 -43
rect 369 -45 372 -43
rect 364 -47 372 -45
rect 374 -40 382 -37
rect 374 -42 377 -40
rect 379 -42 382 -40
rect 374 -44 382 -42
rect 384 -32 392 -30
rect 384 -34 387 -32
rect 389 -34 392 -32
rect 384 -44 392 -34
rect 394 -32 401 -30
rect 394 -34 397 -32
rect 399 -34 401 -32
rect 394 -39 401 -34
rect 407 -37 412 -30
rect 394 -41 397 -39
rect 399 -41 401 -39
rect 394 -44 401 -41
rect 405 -39 412 -37
rect 405 -41 407 -39
rect 409 -41 412 -39
rect 405 -43 412 -41
rect 374 -47 379 -44
rect 364 -50 369 -47
rect 407 -50 412 -43
rect 414 -50 419 -30
rect 421 -36 428 -30
rect 456 -36 463 -30
rect 421 -46 430 -36
rect 421 -48 424 -46
rect 426 -48 430 -46
rect 421 -50 430 -48
rect 432 -39 439 -36
rect 432 -41 435 -39
rect 437 -41 439 -39
rect 432 -43 439 -41
rect 445 -39 452 -36
rect 445 -41 447 -39
rect 449 -41 452 -39
rect 445 -43 452 -41
rect 432 -50 437 -43
rect 447 -50 452 -43
rect 454 -46 463 -36
rect 454 -48 458 -46
rect 460 -48 463 -46
rect 454 -50 463 -48
rect 465 -50 470 -30
rect 472 -37 477 -30
rect 483 -32 490 -30
rect 483 -34 485 -32
rect 487 -34 490 -32
rect 472 -39 479 -37
rect 472 -41 475 -39
rect 477 -41 479 -39
rect 472 -43 479 -41
rect 483 -39 490 -34
rect 483 -41 485 -39
rect 487 -41 490 -39
rect 472 -50 477 -43
rect 483 -44 490 -41
rect 492 -32 500 -30
rect 492 -34 495 -32
rect 497 -34 500 -32
rect 492 -44 500 -34
rect 502 -37 507 -30
rect 534 -36 541 -30
rect 543 -32 551 -30
rect 543 -34 546 -32
rect 548 -34 551 -32
rect 543 -36 551 -34
rect 553 -36 561 -30
rect 502 -40 510 -37
rect 502 -42 505 -40
rect 507 -42 510 -40
rect 502 -44 510 -42
rect 505 -47 510 -44
rect 512 -43 520 -37
rect 512 -45 515 -43
rect 517 -45 520 -43
rect 512 -47 520 -45
rect 515 -50 520 -47
rect 522 -39 529 -37
rect 522 -41 525 -39
rect 527 -41 529 -39
rect 522 -43 529 -41
rect 534 -43 539 -36
rect 555 -39 561 -36
rect 563 -32 570 -30
rect 563 -34 566 -32
rect 568 -34 570 -32
rect 563 -36 570 -34
rect 563 -39 568 -36
rect 584 -37 589 -32
rect 582 -39 589 -37
rect 555 -43 559 -39
rect 522 -50 527 -43
rect 534 -45 540 -43
rect 534 -47 536 -45
rect 538 -47 540 -45
rect 534 -49 540 -47
rect 553 -45 559 -43
rect 582 -41 584 -39
rect 586 -41 589 -39
rect 582 -43 589 -41
rect 591 -43 596 -32
rect 598 -41 609 -32
rect 611 -35 616 -32
rect 611 -37 618 -35
rect 644 -37 649 -30
rect 611 -39 614 -37
rect 616 -39 618 -37
rect 611 -41 618 -39
rect 622 -39 629 -37
rect 622 -41 624 -39
rect 626 -41 629 -39
rect 598 -43 607 -41
rect 553 -47 555 -45
rect 557 -47 559 -45
rect 553 -49 559 -47
rect 600 -49 607 -43
rect 622 -43 629 -41
rect 600 -51 603 -49
rect 605 -51 607 -49
rect 600 -53 607 -51
rect 624 -50 629 -43
rect 631 -43 639 -37
rect 631 -45 634 -43
rect 636 -45 639 -43
rect 631 -47 639 -45
rect 641 -40 649 -37
rect 641 -42 644 -40
rect 646 -42 649 -40
rect 641 -44 649 -42
rect 651 -32 659 -30
rect 651 -34 654 -32
rect 656 -34 659 -32
rect 651 -44 659 -34
rect 661 -32 668 -30
rect 661 -34 664 -32
rect 666 -34 668 -32
rect 661 -39 668 -34
rect 674 -37 679 -30
rect 661 -41 664 -39
rect 666 -41 668 -39
rect 661 -44 668 -41
rect 672 -39 679 -37
rect 672 -41 674 -39
rect 676 -41 679 -39
rect 672 -43 679 -41
rect 641 -47 646 -44
rect 631 -50 636 -47
rect 674 -50 679 -43
rect 681 -50 686 -30
rect 688 -36 695 -30
rect 723 -36 730 -30
rect 688 -46 697 -36
rect 688 -48 691 -46
rect 693 -48 697 -46
rect 688 -50 697 -48
rect 699 -39 706 -36
rect 699 -41 702 -39
rect 704 -41 706 -39
rect 699 -43 706 -41
rect 712 -39 719 -36
rect 712 -41 714 -39
rect 716 -41 719 -39
rect 712 -43 719 -41
rect 699 -50 704 -43
rect 714 -50 719 -43
rect 721 -46 730 -36
rect 721 -48 725 -46
rect 727 -48 730 -46
rect 721 -50 730 -48
rect 732 -50 737 -30
rect 739 -37 744 -30
rect 750 -32 757 -30
rect 750 -34 752 -32
rect 754 -34 757 -32
rect 739 -39 746 -37
rect 739 -41 742 -39
rect 744 -41 746 -39
rect 739 -43 746 -41
rect 750 -39 757 -34
rect 750 -41 752 -39
rect 754 -41 757 -39
rect 739 -50 744 -43
rect 750 -44 757 -41
rect 759 -32 767 -30
rect 759 -34 762 -32
rect 764 -34 767 -32
rect 759 -44 767 -34
rect 769 -37 774 -30
rect 801 -36 808 -30
rect 810 -32 818 -30
rect 810 -34 813 -32
rect 815 -34 818 -32
rect 810 -36 818 -34
rect 820 -36 828 -30
rect 769 -40 777 -37
rect 769 -42 772 -40
rect 774 -42 777 -40
rect 769 -44 777 -42
rect 772 -47 777 -44
rect 779 -43 787 -37
rect 779 -45 782 -43
rect 784 -45 787 -43
rect 779 -47 787 -45
rect 782 -50 787 -47
rect 789 -39 796 -37
rect 789 -41 792 -39
rect 794 -41 796 -39
rect 789 -43 796 -41
rect 801 -43 806 -36
rect 822 -39 828 -36
rect 830 -32 837 -30
rect 830 -34 833 -32
rect 835 -34 837 -32
rect 830 -36 837 -34
rect 830 -39 835 -36
rect 851 -37 856 -32
rect 849 -39 856 -37
rect 822 -43 826 -39
rect 789 -50 794 -43
rect 801 -45 807 -43
rect 801 -47 803 -45
rect 805 -47 807 -45
rect 801 -49 807 -47
rect 820 -45 826 -43
rect 849 -41 851 -39
rect 853 -41 856 -39
rect 849 -43 856 -41
rect 858 -43 863 -32
rect 865 -41 876 -32
rect 878 -35 883 -32
rect 878 -37 885 -35
rect 911 -37 916 -30
rect 878 -39 881 -37
rect 883 -39 885 -37
rect 878 -41 885 -39
rect 889 -39 896 -37
rect 889 -41 891 -39
rect 893 -41 896 -39
rect 865 -43 874 -41
rect 820 -47 822 -45
rect 824 -47 826 -45
rect 820 -49 826 -47
rect 867 -49 874 -43
rect 889 -43 896 -41
rect 867 -51 870 -49
rect 872 -51 874 -49
rect 867 -53 874 -51
rect 891 -50 896 -43
rect 898 -43 906 -37
rect 898 -45 901 -43
rect 903 -45 906 -43
rect 898 -47 906 -45
rect 908 -40 916 -37
rect 908 -42 911 -40
rect 913 -42 916 -40
rect 908 -44 916 -42
rect 918 -32 926 -30
rect 918 -34 921 -32
rect 923 -34 926 -32
rect 918 -44 926 -34
rect 928 -32 935 -30
rect 928 -34 931 -32
rect 933 -34 935 -32
rect 928 -39 935 -34
rect 941 -37 946 -30
rect 928 -41 931 -39
rect 933 -41 935 -39
rect 928 -44 935 -41
rect 939 -39 946 -37
rect 939 -41 941 -39
rect 943 -41 946 -39
rect 939 -43 946 -41
rect 908 -47 913 -44
rect 898 -50 903 -47
rect 941 -50 946 -43
rect 948 -50 953 -30
rect 955 -36 962 -30
rect 990 -36 997 -30
rect 955 -46 964 -36
rect 955 -48 958 -46
rect 960 -48 964 -46
rect 955 -50 964 -48
rect 966 -39 973 -36
rect 966 -41 969 -39
rect 971 -41 973 -39
rect 966 -43 973 -41
rect 979 -39 986 -36
rect 979 -41 981 -39
rect 983 -41 986 -39
rect 979 -43 986 -41
rect 966 -50 971 -43
rect 981 -50 986 -43
rect 988 -46 997 -36
rect 988 -48 992 -46
rect 994 -48 997 -46
rect 988 -50 997 -48
rect 999 -50 1004 -30
rect 1006 -37 1011 -30
rect 1017 -32 1024 -30
rect 1017 -34 1019 -32
rect 1021 -34 1024 -32
rect 1006 -39 1013 -37
rect 1006 -41 1009 -39
rect 1011 -41 1013 -39
rect 1006 -43 1013 -41
rect 1017 -39 1024 -34
rect 1017 -41 1019 -39
rect 1021 -41 1024 -39
rect 1006 -50 1011 -43
rect 1017 -44 1024 -41
rect 1026 -32 1034 -30
rect 1026 -34 1029 -32
rect 1031 -34 1034 -32
rect 1026 -44 1034 -34
rect 1036 -37 1041 -30
rect 1068 -36 1075 -30
rect 1077 -32 1085 -30
rect 1077 -34 1080 -32
rect 1082 -34 1085 -32
rect 1077 -36 1085 -34
rect 1087 -36 1095 -30
rect 1036 -40 1044 -37
rect 1036 -42 1039 -40
rect 1041 -42 1044 -40
rect 1036 -44 1044 -42
rect 1039 -47 1044 -44
rect 1046 -43 1054 -37
rect 1046 -45 1049 -43
rect 1051 -45 1054 -43
rect 1046 -47 1054 -45
rect 1049 -50 1054 -47
rect 1056 -39 1063 -37
rect 1056 -41 1059 -39
rect 1061 -41 1063 -39
rect 1056 -43 1063 -41
rect 1068 -43 1073 -36
rect 1089 -39 1095 -36
rect 1097 -32 1104 -30
rect 1097 -34 1100 -32
rect 1102 -34 1104 -32
rect 1097 -36 1104 -34
rect 1097 -39 1102 -36
rect 1118 -37 1123 -32
rect 1116 -39 1123 -37
rect 1089 -43 1093 -39
rect 1056 -50 1061 -43
rect 1068 -45 1074 -43
rect 1068 -47 1070 -45
rect 1072 -47 1074 -45
rect 1068 -49 1074 -47
rect 1087 -45 1093 -43
rect 1116 -41 1118 -39
rect 1120 -41 1123 -39
rect 1116 -43 1123 -41
rect 1125 -43 1130 -32
rect 1132 -41 1143 -32
rect 1145 -35 1150 -32
rect 1145 -37 1152 -35
rect 1178 -37 1183 -30
rect 1145 -39 1148 -37
rect 1150 -39 1152 -37
rect 1145 -41 1152 -39
rect 1156 -39 1163 -37
rect 1156 -41 1158 -39
rect 1160 -41 1163 -39
rect 1132 -43 1141 -41
rect 1087 -47 1089 -45
rect 1091 -47 1093 -45
rect 1087 -49 1093 -47
rect 1134 -49 1141 -43
rect 1156 -43 1163 -41
rect 1134 -51 1137 -49
rect 1139 -51 1141 -49
rect 1134 -53 1141 -51
rect 1158 -50 1163 -43
rect 1165 -43 1173 -37
rect 1165 -45 1168 -43
rect 1170 -45 1173 -43
rect 1165 -47 1173 -45
rect 1175 -40 1183 -37
rect 1175 -42 1178 -40
rect 1180 -42 1183 -40
rect 1175 -44 1183 -42
rect 1185 -32 1193 -30
rect 1185 -34 1188 -32
rect 1190 -34 1193 -32
rect 1185 -44 1193 -34
rect 1195 -32 1202 -30
rect 1195 -34 1198 -32
rect 1200 -34 1202 -32
rect 1195 -39 1202 -34
rect 1208 -37 1213 -30
rect 1195 -41 1198 -39
rect 1200 -41 1202 -39
rect 1195 -44 1202 -41
rect 1206 -39 1213 -37
rect 1206 -41 1208 -39
rect 1210 -41 1213 -39
rect 1206 -43 1213 -41
rect 1175 -47 1180 -44
rect 1165 -50 1170 -47
rect 1208 -50 1213 -43
rect 1215 -50 1220 -30
rect 1222 -36 1229 -30
rect 1257 -36 1264 -30
rect 1222 -46 1231 -36
rect 1222 -48 1225 -46
rect 1227 -48 1231 -46
rect 1222 -50 1231 -48
rect 1233 -39 1240 -36
rect 1233 -41 1236 -39
rect 1238 -41 1240 -39
rect 1233 -43 1240 -41
rect 1246 -39 1253 -36
rect 1246 -41 1248 -39
rect 1250 -41 1253 -39
rect 1246 -43 1253 -41
rect 1233 -50 1238 -43
rect 1248 -50 1253 -43
rect 1255 -46 1264 -36
rect 1255 -48 1259 -46
rect 1261 -48 1264 -46
rect 1255 -50 1264 -48
rect 1266 -50 1271 -30
rect 1273 -37 1278 -30
rect 1284 -32 1291 -30
rect 1284 -34 1286 -32
rect 1288 -34 1291 -32
rect 1273 -39 1280 -37
rect 1273 -41 1276 -39
rect 1278 -41 1280 -39
rect 1273 -43 1280 -41
rect 1284 -39 1291 -34
rect 1284 -41 1286 -39
rect 1288 -41 1291 -39
rect 1273 -50 1278 -43
rect 1284 -44 1291 -41
rect 1293 -32 1301 -30
rect 1293 -34 1296 -32
rect 1298 -34 1301 -32
rect 1293 -44 1301 -34
rect 1303 -37 1308 -30
rect 1335 -36 1342 -30
rect 1344 -32 1352 -30
rect 1344 -34 1347 -32
rect 1349 -34 1352 -32
rect 1344 -36 1352 -34
rect 1354 -36 1362 -30
rect 1303 -40 1311 -37
rect 1303 -42 1306 -40
rect 1308 -42 1311 -40
rect 1303 -44 1311 -42
rect 1306 -47 1311 -44
rect 1313 -43 1321 -37
rect 1313 -45 1316 -43
rect 1318 -45 1321 -43
rect 1313 -47 1321 -45
rect 1316 -50 1321 -47
rect 1323 -39 1330 -37
rect 1323 -41 1326 -39
rect 1328 -41 1330 -39
rect 1323 -43 1330 -41
rect 1335 -43 1340 -36
rect 1356 -39 1362 -36
rect 1364 -32 1371 -30
rect 1364 -34 1367 -32
rect 1369 -34 1371 -32
rect 1364 -36 1371 -34
rect 1364 -39 1369 -36
rect 1385 -37 1390 -32
rect 1383 -39 1390 -37
rect 1356 -43 1360 -39
rect 1323 -50 1328 -43
rect 1335 -45 1341 -43
rect 1335 -47 1337 -45
rect 1339 -47 1341 -45
rect 1335 -49 1341 -47
rect 1354 -45 1360 -43
rect 1383 -41 1385 -39
rect 1387 -41 1390 -39
rect 1383 -43 1390 -41
rect 1392 -43 1397 -32
rect 1399 -41 1410 -32
rect 1412 -35 1417 -32
rect 1412 -37 1419 -35
rect 1445 -37 1450 -30
rect 1412 -39 1415 -37
rect 1417 -39 1419 -37
rect 1412 -41 1419 -39
rect 1423 -39 1430 -37
rect 1423 -41 1425 -39
rect 1427 -41 1430 -39
rect 1399 -43 1408 -41
rect 1354 -47 1356 -45
rect 1358 -47 1360 -45
rect 1354 -49 1360 -47
rect 1401 -49 1408 -43
rect 1423 -43 1430 -41
rect 1401 -51 1404 -49
rect 1406 -51 1408 -49
rect 1401 -53 1408 -51
rect 1425 -50 1430 -43
rect 1432 -43 1440 -37
rect 1432 -45 1435 -43
rect 1437 -45 1440 -43
rect 1432 -47 1440 -45
rect 1442 -40 1450 -37
rect 1442 -42 1445 -40
rect 1447 -42 1450 -40
rect 1442 -44 1450 -42
rect 1452 -32 1460 -30
rect 1452 -34 1455 -32
rect 1457 -34 1460 -32
rect 1452 -44 1460 -34
rect 1462 -32 1469 -30
rect 1462 -34 1465 -32
rect 1467 -34 1469 -32
rect 1462 -39 1469 -34
rect 1475 -37 1480 -30
rect 1462 -41 1465 -39
rect 1467 -41 1469 -39
rect 1462 -44 1469 -41
rect 1473 -39 1480 -37
rect 1473 -41 1475 -39
rect 1477 -41 1480 -39
rect 1473 -43 1480 -41
rect 1442 -47 1447 -44
rect 1432 -50 1437 -47
rect 1475 -50 1480 -43
rect 1482 -50 1487 -30
rect 1489 -36 1496 -30
rect 1524 -36 1531 -30
rect 1489 -46 1498 -36
rect 1489 -48 1492 -46
rect 1494 -48 1498 -46
rect 1489 -50 1498 -48
rect 1500 -39 1507 -36
rect 1500 -41 1503 -39
rect 1505 -41 1507 -39
rect 1500 -43 1507 -41
rect 1513 -39 1520 -36
rect 1513 -41 1515 -39
rect 1517 -41 1520 -39
rect 1513 -43 1520 -41
rect 1500 -50 1505 -43
rect 1515 -50 1520 -43
rect 1522 -46 1531 -36
rect 1522 -48 1526 -46
rect 1528 -48 1531 -46
rect 1522 -50 1531 -48
rect 1533 -50 1538 -30
rect 1540 -37 1545 -30
rect 1551 -32 1558 -30
rect 1551 -34 1553 -32
rect 1555 -34 1558 -32
rect 1540 -39 1547 -37
rect 1540 -41 1543 -39
rect 1545 -41 1547 -39
rect 1540 -43 1547 -41
rect 1551 -39 1558 -34
rect 1551 -41 1553 -39
rect 1555 -41 1558 -39
rect 1540 -50 1545 -43
rect 1551 -44 1558 -41
rect 1560 -32 1568 -30
rect 1560 -34 1563 -32
rect 1565 -34 1568 -32
rect 1560 -44 1568 -34
rect 1570 -37 1575 -30
rect 1602 -36 1609 -30
rect 1611 -32 1619 -30
rect 1611 -34 1614 -32
rect 1616 -34 1619 -32
rect 1611 -36 1619 -34
rect 1621 -36 1629 -30
rect 1570 -40 1578 -37
rect 1570 -42 1573 -40
rect 1575 -42 1578 -40
rect 1570 -44 1578 -42
rect 1573 -47 1578 -44
rect 1580 -43 1588 -37
rect 1580 -45 1583 -43
rect 1585 -45 1588 -43
rect 1580 -47 1588 -45
rect 1583 -50 1588 -47
rect 1590 -39 1597 -37
rect 1590 -41 1593 -39
rect 1595 -41 1597 -39
rect 1590 -43 1597 -41
rect 1602 -43 1607 -36
rect 1623 -39 1629 -36
rect 1631 -32 1638 -30
rect 1631 -34 1634 -32
rect 1636 -34 1638 -32
rect 1631 -36 1638 -34
rect 1631 -39 1636 -36
rect 1652 -37 1657 -32
rect 1650 -39 1657 -37
rect 1623 -43 1627 -39
rect 1590 -50 1595 -43
rect 1602 -45 1608 -43
rect 1602 -47 1604 -45
rect 1606 -47 1608 -45
rect 1602 -49 1608 -47
rect 1621 -45 1627 -43
rect 1650 -41 1652 -39
rect 1654 -41 1657 -39
rect 1650 -43 1657 -41
rect 1659 -43 1664 -32
rect 1666 -41 1677 -32
rect 1679 -35 1684 -32
rect 1679 -37 1686 -35
rect 1712 -37 1717 -30
rect 1679 -39 1682 -37
rect 1684 -39 1686 -37
rect 1679 -41 1686 -39
rect 1690 -39 1697 -37
rect 1690 -41 1692 -39
rect 1694 -41 1697 -39
rect 1666 -43 1675 -41
rect 1621 -47 1623 -45
rect 1625 -47 1627 -45
rect 1621 -49 1627 -47
rect 1668 -49 1675 -43
rect 1690 -43 1697 -41
rect 1668 -51 1671 -49
rect 1673 -51 1675 -49
rect 1668 -53 1675 -51
rect 1692 -50 1697 -43
rect 1699 -43 1707 -37
rect 1699 -45 1702 -43
rect 1704 -45 1707 -43
rect 1699 -47 1707 -45
rect 1709 -40 1717 -37
rect 1709 -42 1712 -40
rect 1714 -42 1717 -40
rect 1709 -44 1717 -42
rect 1719 -32 1727 -30
rect 1719 -34 1722 -32
rect 1724 -34 1727 -32
rect 1719 -44 1727 -34
rect 1729 -32 1736 -30
rect 1729 -34 1732 -32
rect 1734 -34 1736 -32
rect 1729 -39 1736 -34
rect 1742 -37 1747 -30
rect 1729 -41 1732 -39
rect 1734 -41 1736 -39
rect 1729 -44 1736 -41
rect 1740 -39 1747 -37
rect 1740 -41 1742 -39
rect 1744 -41 1747 -39
rect 1740 -43 1747 -41
rect 1709 -47 1714 -44
rect 1699 -50 1704 -47
rect 1742 -50 1747 -43
rect 1749 -50 1754 -30
rect 1756 -36 1763 -30
rect 1791 -36 1798 -30
rect 1756 -46 1765 -36
rect 1756 -48 1759 -46
rect 1761 -48 1765 -46
rect 1756 -50 1765 -48
rect 1767 -39 1774 -36
rect 1767 -41 1770 -39
rect 1772 -41 1774 -39
rect 1767 -43 1774 -41
rect 1780 -39 1787 -36
rect 1780 -41 1782 -39
rect 1784 -41 1787 -39
rect 1780 -43 1787 -41
rect 1767 -50 1772 -43
rect 1782 -50 1787 -43
rect 1789 -46 1798 -36
rect 1789 -48 1793 -46
rect 1795 -48 1798 -46
rect 1789 -50 1798 -48
rect 1800 -50 1805 -30
rect 1807 -37 1812 -30
rect 1818 -32 1825 -30
rect 1818 -34 1820 -32
rect 1822 -34 1825 -32
rect 1807 -39 1814 -37
rect 1807 -41 1810 -39
rect 1812 -41 1814 -39
rect 1807 -43 1814 -41
rect 1818 -39 1825 -34
rect 1818 -41 1820 -39
rect 1822 -41 1825 -39
rect 1807 -50 1812 -43
rect 1818 -44 1825 -41
rect 1827 -32 1835 -30
rect 1827 -34 1830 -32
rect 1832 -34 1835 -32
rect 1827 -44 1835 -34
rect 1837 -37 1842 -30
rect 1869 -36 1876 -30
rect 1878 -32 1886 -30
rect 1878 -34 1881 -32
rect 1883 -34 1886 -32
rect 1878 -36 1886 -34
rect 1888 -36 1896 -30
rect 1837 -40 1845 -37
rect 1837 -42 1840 -40
rect 1842 -42 1845 -40
rect 1837 -44 1845 -42
rect 1840 -47 1845 -44
rect 1847 -43 1855 -37
rect 1847 -45 1850 -43
rect 1852 -45 1855 -43
rect 1847 -47 1855 -45
rect 1850 -50 1855 -47
rect 1857 -39 1864 -37
rect 1857 -41 1860 -39
rect 1862 -41 1864 -39
rect 1857 -43 1864 -41
rect 1869 -43 1874 -36
rect 1890 -39 1896 -36
rect 1898 -32 1905 -30
rect 1898 -34 1901 -32
rect 1903 -34 1905 -32
rect 1898 -36 1905 -34
rect 1912 -32 1919 -30
rect 1912 -34 1914 -32
rect 1916 -34 1919 -32
rect 1912 -36 1919 -34
rect 1898 -39 1903 -36
rect 1914 -39 1919 -36
rect 1921 -35 1926 -30
rect 1921 -39 1935 -35
rect 1890 -43 1894 -39
rect 1857 -50 1862 -43
rect 1869 -45 1875 -43
rect 1869 -47 1871 -45
rect 1873 -47 1875 -45
rect 1869 -49 1875 -47
rect 1888 -45 1894 -43
rect 1926 -40 1935 -39
rect 1926 -42 1928 -40
rect 1930 -42 1935 -40
rect 1926 -44 1935 -42
rect 1937 -37 1945 -35
rect 1937 -39 1940 -37
rect 1942 -39 1945 -37
rect 1937 -44 1945 -39
rect 1947 -39 1955 -35
rect 1947 -41 1950 -39
rect 1952 -41 1955 -39
rect 1947 -44 1955 -41
rect 1888 -47 1890 -45
rect 1892 -47 1894 -45
rect 1888 -49 1894 -47
rect 1950 -47 1955 -44
rect 1957 -47 1962 -35
rect 1964 -47 1972 -35
rect 1998 -37 2003 -30
rect 1976 -39 1983 -37
rect 1976 -41 1978 -39
rect 1980 -41 1983 -39
rect 1976 -43 1983 -41
rect 1966 -49 1972 -47
rect 1966 -51 1968 -49
rect 1970 -51 1972 -49
rect 1978 -50 1983 -43
rect 1985 -43 1993 -37
rect 1985 -45 1988 -43
rect 1990 -45 1993 -43
rect 1985 -47 1993 -45
rect 1995 -40 2003 -37
rect 1995 -42 1998 -40
rect 2000 -42 2003 -40
rect 1995 -44 2003 -42
rect 2005 -32 2013 -30
rect 2005 -34 2008 -32
rect 2010 -34 2013 -32
rect 2005 -44 2013 -34
rect 2015 -32 2022 -30
rect 2015 -34 2018 -32
rect 2020 -34 2022 -32
rect 2015 -39 2022 -34
rect 2028 -37 2033 -30
rect 2015 -41 2018 -39
rect 2020 -41 2022 -39
rect 2015 -44 2022 -41
rect 2026 -39 2033 -37
rect 2026 -41 2028 -39
rect 2030 -41 2033 -39
rect 2026 -43 2033 -41
rect 1995 -47 2000 -44
rect 1985 -50 1990 -47
rect 1966 -53 1972 -51
rect 2028 -50 2033 -43
rect 2035 -50 2040 -30
rect 2042 -36 2049 -30
rect 2077 -36 2084 -30
rect 2042 -46 2051 -36
rect 2042 -48 2045 -46
rect 2047 -48 2051 -46
rect 2042 -50 2051 -48
rect 2053 -39 2060 -36
rect 2053 -41 2056 -39
rect 2058 -41 2060 -39
rect 2053 -43 2060 -41
rect 2066 -39 2073 -36
rect 2066 -41 2068 -39
rect 2070 -41 2073 -39
rect 2066 -43 2073 -41
rect 2053 -50 2058 -43
rect 2068 -50 2073 -43
rect 2075 -46 2084 -36
rect 2075 -48 2079 -46
rect 2081 -48 2084 -46
rect 2075 -50 2084 -48
rect 2086 -50 2091 -30
rect 2093 -37 2098 -30
rect 2104 -32 2111 -30
rect 2104 -34 2106 -32
rect 2108 -34 2111 -32
rect 2093 -39 2100 -37
rect 2093 -41 2096 -39
rect 2098 -41 2100 -39
rect 2093 -43 2100 -41
rect 2104 -39 2111 -34
rect 2104 -41 2106 -39
rect 2108 -41 2111 -39
rect 2093 -50 2098 -43
rect 2104 -44 2111 -41
rect 2113 -32 2121 -30
rect 2113 -34 2116 -32
rect 2118 -34 2121 -32
rect 2113 -44 2121 -34
rect 2123 -37 2128 -30
rect 2155 -36 2162 -30
rect 2164 -32 2172 -30
rect 2164 -34 2167 -32
rect 2169 -34 2172 -32
rect 2164 -36 2172 -34
rect 2174 -36 2182 -30
rect 2123 -40 2131 -37
rect 2123 -42 2126 -40
rect 2128 -42 2131 -40
rect 2123 -44 2131 -42
rect 2126 -47 2131 -44
rect 2133 -43 2141 -37
rect 2133 -45 2136 -43
rect 2138 -45 2141 -43
rect 2133 -47 2141 -45
rect 2136 -50 2141 -47
rect 2143 -39 2150 -37
rect 2143 -41 2146 -39
rect 2148 -41 2150 -39
rect 2143 -43 2150 -41
rect 2155 -43 2160 -36
rect 2176 -39 2182 -36
rect 2184 -32 2191 -30
rect 2184 -34 2187 -32
rect 2189 -34 2191 -32
rect 2184 -36 2191 -34
rect 2245 -36 2250 -35
rect 2184 -39 2189 -36
rect 2199 -38 2206 -36
rect 2176 -43 2180 -39
rect 2143 -50 2148 -43
rect 2155 -45 2161 -43
rect 2155 -47 2157 -45
rect 2159 -47 2161 -45
rect 2155 -49 2161 -47
rect 2174 -45 2180 -43
rect 2199 -40 2201 -38
rect 2203 -40 2206 -38
rect 2199 -42 2206 -40
rect 2208 -38 2216 -36
rect 2208 -40 2211 -38
rect 2213 -40 2216 -38
rect 2208 -42 2216 -40
rect 2174 -47 2176 -45
rect 2178 -47 2180 -45
rect 2174 -49 2180 -47
rect 2210 -44 2216 -42
rect 2218 -44 2223 -36
rect 2225 -40 2233 -36
rect 2225 -42 2228 -40
rect 2230 -42 2233 -40
rect 2225 -44 2233 -42
rect 2235 -44 2240 -36
rect 2242 -40 2250 -36
rect 2242 -42 2245 -40
rect 2247 -42 2250 -40
rect 2242 -44 2250 -42
rect 2252 -37 2259 -35
rect 2313 -36 2318 -35
rect 2252 -39 2255 -37
rect 2257 -39 2259 -37
rect 2252 -41 2259 -39
rect 2267 -38 2274 -36
rect 2267 -40 2269 -38
rect 2271 -40 2274 -38
rect 2252 -44 2257 -41
rect 2267 -42 2274 -40
rect 2276 -38 2284 -36
rect 2276 -40 2279 -38
rect 2281 -40 2284 -38
rect 2276 -42 2284 -40
rect 2278 -44 2284 -42
rect 2286 -44 2291 -36
rect 2293 -40 2301 -36
rect 2293 -42 2296 -40
rect 2298 -42 2301 -40
rect 2293 -44 2301 -42
rect 2303 -44 2308 -36
rect 2310 -40 2318 -36
rect 2310 -42 2313 -40
rect 2315 -42 2318 -40
rect 2310 -44 2318 -42
rect 2320 -37 2327 -35
rect 2320 -39 2323 -37
rect 2325 -39 2327 -37
rect 2320 -41 2327 -39
rect 2320 -44 2325 -41
rect 26 -61 33 -59
rect 26 -63 29 -61
rect 31 -63 33 -61
rect 26 -69 33 -63
rect 66 -61 73 -59
rect 66 -63 69 -61
rect 71 -63 73 -61
rect 8 -71 15 -69
rect 8 -73 10 -71
rect 12 -73 15 -71
rect 8 -75 15 -73
rect 10 -80 15 -75
rect 17 -80 22 -69
rect 24 -71 33 -69
rect 66 -69 73 -63
rect 48 -71 55 -69
rect 24 -80 35 -71
rect 37 -73 44 -71
rect 37 -75 40 -73
rect 42 -75 44 -73
rect 48 -73 50 -71
rect 52 -73 55 -71
rect 48 -75 55 -73
rect 37 -77 44 -75
rect 37 -80 42 -77
rect 50 -80 55 -75
rect 57 -80 62 -69
rect 64 -71 73 -69
rect 90 -69 95 -62
rect 88 -71 95 -69
rect 64 -80 75 -71
rect 77 -73 84 -71
rect 77 -75 80 -73
rect 82 -75 84 -73
rect 88 -73 90 -71
rect 92 -73 95 -71
rect 88 -75 95 -73
rect 97 -65 102 -62
rect 97 -67 105 -65
rect 97 -69 100 -67
rect 102 -69 105 -67
rect 97 -75 105 -69
rect 107 -68 112 -65
rect 107 -70 115 -68
rect 107 -72 110 -70
rect 112 -72 115 -70
rect 107 -75 115 -72
rect 77 -77 84 -75
rect 77 -80 82 -77
rect 110 -82 115 -75
rect 117 -78 125 -68
rect 117 -80 120 -78
rect 122 -80 125 -78
rect 117 -82 125 -80
rect 127 -71 134 -68
rect 140 -69 145 -62
rect 127 -73 130 -71
rect 132 -73 134 -71
rect 127 -78 134 -73
rect 138 -71 145 -69
rect 138 -73 140 -71
rect 142 -73 145 -71
rect 138 -75 145 -73
rect 127 -80 130 -78
rect 132 -80 134 -78
rect 127 -82 134 -80
rect 140 -82 145 -75
rect 147 -82 152 -62
rect 154 -64 163 -62
rect 154 -66 157 -64
rect 159 -66 163 -64
rect 154 -76 163 -66
rect 165 -69 170 -62
rect 180 -69 185 -62
rect 165 -71 172 -69
rect 165 -73 168 -71
rect 170 -73 172 -71
rect 165 -76 172 -73
rect 178 -71 185 -69
rect 178 -73 180 -71
rect 182 -73 185 -71
rect 178 -76 185 -73
rect 187 -64 196 -62
rect 187 -66 191 -64
rect 193 -66 196 -64
rect 187 -76 196 -66
rect 154 -82 161 -76
rect 189 -82 196 -76
rect 198 -82 203 -62
rect 205 -69 210 -62
rect 248 -65 253 -62
rect 238 -68 243 -65
rect 205 -71 212 -69
rect 205 -73 208 -71
rect 210 -73 212 -71
rect 205 -75 212 -73
rect 216 -71 223 -68
rect 216 -73 218 -71
rect 220 -73 223 -71
rect 205 -82 210 -75
rect 216 -78 223 -73
rect 216 -80 218 -78
rect 220 -80 223 -78
rect 216 -82 223 -80
rect 225 -78 233 -68
rect 225 -80 228 -78
rect 230 -80 233 -78
rect 225 -82 233 -80
rect 235 -70 243 -68
rect 235 -72 238 -70
rect 240 -72 243 -70
rect 235 -75 243 -72
rect 245 -67 253 -65
rect 245 -69 248 -67
rect 250 -69 253 -67
rect 245 -75 253 -69
rect 255 -69 260 -62
rect 267 -65 273 -63
rect 267 -67 269 -65
rect 271 -67 273 -65
rect 267 -69 273 -67
rect 286 -65 292 -63
rect 333 -61 340 -59
rect 333 -63 336 -61
rect 338 -63 340 -61
rect 286 -67 288 -65
rect 290 -67 292 -65
rect 286 -69 292 -67
rect 255 -71 262 -69
rect 255 -73 258 -71
rect 260 -73 262 -71
rect 255 -75 262 -73
rect 235 -82 240 -75
rect 267 -76 272 -69
rect 288 -73 292 -69
rect 333 -69 340 -63
rect 315 -71 322 -69
rect 315 -73 317 -71
rect 319 -73 322 -71
rect 288 -76 294 -73
rect 267 -82 274 -76
rect 276 -78 284 -76
rect 276 -80 279 -78
rect 281 -80 284 -78
rect 276 -82 284 -80
rect 286 -82 294 -76
rect 296 -76 301 -73
rect 315 -75 322 -73
rect 296 -78 303 -76
rect 296 -80 299 -78
rect 301 -80 303 -78
rect 317 -80 322 -75
rect 324 -80 329 -69
rect 331 -71 340 -69
rect 357 -69 362 -62
rect 355 -71 362 -69
rect 331 -80 342 -71
rect 344 -73 351 -71
rect 344 -75 347 -73
rect 349 -75 351 -73
rect 355 -73 357 -71
rect 359 -73 362 -71
rect 355 -75 362 -73
rect 364 -65 369 -62
rect 364 -67 372 -65
rect 364 -69 367 -67
rect 369 -69 372 -67
rect 364 -75 372 -69
rect 374 -68 379 -65
rect 374 -70 382 -68
rect 374 -72 377 -70
rect 379 -72 382 -70
rect 374 -75 382 -72
rect 344 -77 351 -75
rect 344 -80 349 -77
rect 296 -82 303 -80
rect 377 -82 382 -75
rect 384 -78 392 -68
rect 384 -80 387 -78
rect 389 -80 392 -78
rect 384 -82 392 -80
rect 394 -71 401 -68
rect 407 -69 412 -62
rect 394 -73 397 -71
rect 399 -73 401 -71
rect 394 -78 401 -73
rect 405 -71 412 -69
rect 405 -73 407 -71
rect 409 -73 412 -71
rect 405 -75 412 -73
rect 394 -80 397 -78
rect 399 -80 401 -78
rect 394 -82 401 -80
rect 407 -82 412 -75
rect 414 -82 419 -62
rect 421 -64 430 -62
rect 421 -66 424 -64
rect 426 -66 430 -64
rect 421 -76 430 -66
rect 432 -69 437 -62
rect 447 -69 452 -62
rect 432 -71 439 -69
rect 432 -73 435 -71
rect 437 -73 439 -71
rect 432 -76 439 -73
rect 445 -71 452 -69
rect 445 -73 447 -71
rect 449 -73 452 -71
rect 445 -76 452 -73
rect 454 -64 463 -62
rect 454 -66 458 -64
rect 460 -66 463 -64
rect 454 -76 463 -66
rect 421 -82 428 -76
rect 456 -82 463 -76
rect 465 -82 470 -62
rect 472 -69 477 -62
rect 515 -65 520 -62
rect 505 -68 510 -65
rect 472 -71 479 -69
rect 472 -73 475 -71
rect 477 -73 479 -71
rect 472 -75 479 -73
rect 483 -71 490 -68
rect 483 -73 485 -71
rect 487 -73 490 -71
rect 472 -82 477 -75
rect 483 -78 490 -73
rect 483 -80 485 -78
rect 487 -80 490 -78
rect 483 -82 490 -80
rect 492 -78 500 -68
rect 492 -80 495 -78
rect 497 -80 500 -78
rect 492 -82 500 -80
rect 502 -70 510 -68
rect 502 -72 505 -70
rect 507 -72 510 -70
rect 502 -75 510 -72
rect 512 -67 520 -65
rect 512 -69 515 -67
rect 517 -69 520 -67
rect 512 -75 520 -69
rect 522 -69 527 -62
rect 534 -65 540 -63
rect 534 -67 536 -65
rect 538 -67 540 -65
rect 534 -69 540 -67
rect 553 -65 559 -63
rect 600 -61 607 -59
rect 600 -63 603 -61
rect 605 -63 607 -61
rect 553 -67 555 -65
rect 557 -67 559 -65
rect 553 -69 559 -67
rect 522 -71 529 -69
rect 522 -73 525 -71
rect 527 -73 529 -71
rect 522 -75 529 -73
rect 502 -82 507 -75
rect 534 -76 539 -69
rect 555 -73 559 -69
rect 600 -69 607 -63
rect 582 -71 589 -69
rect 582 -73 584 -71
rect 586 -73 589 -71
rect 555 -76 561 -73
rect 534 -82 541 -76
rect 543 -78 551 -76
rect 543 -80 546 -78
rect 548 -80 551 -78
rect 543 -82 551 -80
rect 553 -82 561 -76
rect 563 -76 568 -73
rect 582 -75 589 -73
rect 563 -78 570 -76
rect 563 -80 566 -78
rect 568 -80 570 -78
rect 584 -80 589 -75
rect 591 -80 596 -69
rect 598 -71 607 -69
rect 624 -69 629 -62
rect 622 -71 629 -69
rect 598 -80 609 -71
rect 611 -73 618 -71
rect 611 -75 614 -73
rect 616 -75 618 -73
rect 622 -73 624 -71
rect 626 -73 629 -71
rect 622 -75 629 -73
rect 631 -65 636 -62
rect 631 -67 639 -65
rect 631 -69 634 -67
rect 636 -69 639 -67
rect 631 -75 639 -69
rect 641 -68 646 -65
rect 641 -70 649 -68
rect 641 -72 644 -70
rect 646 -72 649 -70
rect 641 -75 649 -72
rect 611 -77 618 -75
rect 611 -80 616 -77
rect 563 -82 570 -80
rect 644 -82 649 -75
rect 651 -78 659 -68
rect 651 -80 654 -78
rect 656 -80 659 -78
rect 651 -82 659 -80
rect 661 -71 668 -68
rect 674 -69 679 -62
rect 661 -73 664 -71
rect 666 -73 668 -71
rect 661 -78 668 -73
rect 672 -71 679 -69
rect 672 -73 674 -71
rect 676 -73 679 -71
rect 672 -75 679 -73
rect 661 -80 664 -78
rect 666 -80 668 -78
rect 661 -82 668 -80
rect 674 -82 679 -75
rect 681 -82 686 -62
rect 688 -64 697 -62
rect 688 -66 691 -64
rect 693 -66 697 -64
rect 688 -76 697 -66
rect 699 -69 704 -62
rect 714 -69 719 -62
rect 699 -71 706 -69
rect 699 -73 702 -71
rect 704 -73 706 -71
rect 699 -76 706 -73
rect 712 -71 719 -69
rect 712 -73 714 -71
rect 716 -73 719 -71
rect 712 -76 719 -73
rect 721 -64 730 -62
rect 721 -66 725 -64
rect 727 -66 730 -64
rect 721 -76 730 -66
rect 688 -82 695 -76
rect 723 -82 730 -76
rect 732 -82 737 -62
rect 739 -69 744 -62
rect 782 -65 787 -62
rect 772 -68 777 -65
rect 739 -71 746 -69
rect 739 -73 742 -71
rect 744 -73 746 -71
rect 739 -75 746 -73
rect 750 -71 757 -68
rect 750 -73 752 -71
rect 754 -73 757 -71
rect 739 -82 744 -75
rect 750 -78 757 -73
rect 750 -80 752 -78
rect 754 -80 757 -78
rect 750 -82 757 -80
rect 759 -78 767 -68
rect 759 -80 762 -78
rect 764 -80 767 -78
rect 759 -82 767 -80
rect 769 -70 777 -68
rect 769 -72 772 -70
rect 774 -72 777 -70
rect 769 -75 777 -72
rect 779 -67 787 -65
rect 779 -69 782 -67
rect 784 -69 787 -67
rect 779 -75 787 -69
rect 789 -69 794 -62
rect 801 -65 807 -63
rect 801 -67 803 -65
rect 805 -67 807 -65
rect 801 -69 807 -67
rect 820 -65 826 -63
rect 867 -61 874 -59
rect 867 -63 870 -61
rect 872 -63 874 -61
rect 820 -67 822 -65
rect 824 -67 826 -65
rect 820 -69 826 -67
rect 789 -71 796 -69
rect 789 -73 792 -71
rect 794 -73 796 -71
rect 789 -75 796 -73
rect 769 -82 774 -75
rect 801 -76 806 -69
rect 822 -73 826 -69
rect 867 -69 874 -63
rect 849 -71 856 -69
rect 849 -73 851 -71
rect 853 -73 856 -71
rect 822 -76 828 -73
rect 801 -82 808 -76
rect 810 -78 818 -76
rect 810 -80 813 -78
rect 815 -80 818 -78
rect 810 -82 818 -80
rect 820 -82 828 -76
rect 830 -76 835 -73
rect 849 -75 856 -73
rect 830 -78 837 -76
rect 830 -80 833 -78
rect 835 -80 837 -78
rect 851 -80 856 -75
rect 858 -80 863 -69
rect 865 -71 874 -69
rect 891 -69 896 -62
rect 889 -71 896 -69
rect 865 -80 876 -71
rect 878 -73 885 -71
rect 878 -75 881 -73
rect 883 -75 885 -73
rect 889 -73 891 -71
rect 893 -73 896 -71
rect 889 -75 896 -73
rect 898 -65 903 -62
rect 898 -67 906 -65
rect 898 -69 901 -67
rect 903 -69 906 -67
rect 898 -75 906 -69
rect 908 -68 913 -65
rect 908 -70 916 -68
rect 908 -72 911 -70
rect 913 -72 916 -70
rect 908 -75 916 -72
rect 878 -77 885 -75
rect 878 -80 883 -77
rect 830 -82 837 -80
rect 911 -82 916 -75
rect 918 -78 926 -68
rect 918 -80 921 -78
rect 923 -80 926 -78
rect 918 -82 926 -80
rect 928 -71 935 -68
rect 941 -69 946 -62
rect 928 -73 931 -71
rect 933 -73 935 -71
rect 928 -78 935 -73
rect 939 -71 946 -69
rect 939 -73 941 -71
rect 943 -73 946 -71
rect 939 -75 946 -73
rect 928 -80 931 -78
rect 933 -80 935 -78
rect 928 -82 935 -80
rect 941 -82 946 -75
rect 948 -82 953 -62
rect 955 -64 964 -62
rect 955 -66 958 -64
rect 960 -66 964 -64
rect 955 -76 964 -66
rect 966 -69 971 -62
rect 981 -69 986 -62
rect 966 -71 973 -69
rect 966 -73 969 -71
rect 971 -73 973 -71
rect 966 -76 973 -73
rect 979 -71 986 -69
rect 979 -73 981 -71
rect 983 -73 986 -71
rect 979 -76 986 -73
rect 988 -64 997 -62
rect 988 -66 992 -64
rect 994 -66 997 -64
rect 988 -76 997 -66
rect 955 -82 962 -76
rect 990 -82 997 -76
rect 999 -82 1004 -62
rect 1006 -69 1011 -62
rect 1049 -65 1054 -62
rect 1039 -68 1044 -65
rect 1006 -71 1013 -69
rect 1006 -73 1009 -71
rect 1011 -73 1013 -71
rect 1006 -75 1013 -73
rect 1017 -71 1024 -68
rect 1017 -73 1019 -71
rect 1021 -73 1024 -71
rect 1006 -82 1011 -75
rect 1017 -78 1024 -73
rect 1017 -80 1019 -78
rect 1021 -80 1024 -78
rect 1017 -82 1024 -80
rect 1026 -78 1034 -68
rect 1026 -80 1029 -78
rect 1031 -80 1034 -78
rect 1026 -82 1034 -80
rect 1036 -70 1044 -68
rect 1036 -72 1039 -70
rect 1041 -72 1044 -70
rect 1036 -75 1044 -72
rect 1046 -67 1054 -65
rect 1046 -69 1049 -67
rect 1051 -69 1054 -67
rect 1046 -75 1054 -69
rect 1056 -69 1061 -62
rect 1068 -65 1074 -63
rect 1068 -67 1070 -65
rect 1072 -67 1074 -65
rect 1068 -69 1074 -67
rect 1087 -65 1093 -63
rect 1134 -61 1141 -59
rect 1134 -63 1137 -61
rect 1139 -63 1141 -61
rect 1087 -67 1089 -65
rect 1091 -67 1093 -65
rect 1087 -69 1093 -67
rect 1056 -71 1063 -69
rect 1056 -73 1059 -71
rect 1061 -73 1063 -71
rect 1056 -75 1063 -73
rect 1036 -82 1041 -75
rect 1068 -76 1073 -69
rect 1089 -73 1093 -69
rect 1134 -69 1141 -63
rect 1116 -71 1123 -69
rect 1116 -73 1118 -71
rect 1120 -73 1123 -71
rect 1089 -76 1095 -73
rect 1068 -82 1075 -76
rect 1077 -78 1085 -76
rect 1077 -80 1080 -78
rect 1082 -80 1085 -78
rect 1077 -82 1085 -80
rect 1087 -82 1095 -76
rect 1097 -76 1102 -73
rect 1116 -75 1123 -73
rect 1097 -78 1104 -76
rect 1097 -80 1100 -78
rect 1102 -80 1104 -78
rect 1118 -80 1123 -75
rect 1125 -80 1130 -69
rect 1132 -71 1141 -69
rect 1158 -69 1163 -62
rect 1156 -71 1163 -69
rect 1132 -80 1143 -71
rect 1145 -73 1152 -71
rect 1145 -75 1148 -73
rect 1150 -75 1152 -73
rect 1156 -73 1158 -71
rect 1160 -73 1163 -71
rect 1156 -75 1163 -73
rect 1165 -65 1170 -62
rect 1165 -67 1173 -65
rect 1165 -69 1168 -67
rect 1170 -69 1173 -67
rect 1165 -75 1173 -69
rect 1175 -68 1180 -65
rect 1175 -70 1183 -68
rect 1175 -72 1178 -70
rect 1180 -72 1183 -70
rect 1175 -75 1183 -72
rect 1145 -77 1152 -75
rect 1145 -80 1150 -77
rect 1097 -82 1104 -80
rect 1178 -82 1183 -75
rect 1185 -78 1193 -68
rect 1185 -80 1188 -78
rect 1190 -80 1193 -78
rect 1185 -82 1193 -80
rect 1195 -71 1202 -68
rect 1208 -69 1213 -62
rect 1195 -73 1198 -71
rect 1200 -73 1202 -71
rect 1195 -78 1202 -73
rect 1206 -71 1213 -69
rect 1206 -73 1208 -71
rect 1210 -73 1213 -71
rect 1206 -75 1213 -73
rect 1195 -80 1198 -78
rect 1200 -80 1202 -78
rect 1195 -82 1202 -80
rect 1208 -82 1213 -75
rect 1215 -82 1220 -62
rect 1222 -64 1231 -62
rect 1222 -66 1225 -64
rect 1227 -66 1231 -64
rect 1222 -76 1231 -66
rect 1233 -69 1238 -62
rect 1248 -69 1253 -62
rect 1233 -71 1240 -69
rect 1233 -73 1236 -71
rect 1238 -73 1240 -71
rect 1233 -76 1240 -73
rect 1246 -71 1253 -69
rect 1246 -73 1248 -71
rect 1250 -73 1253 -71
rect 1246 -76 1253 -73
rect 1255 -64 1264 -62
rect 1255 -66 1259 -64
rect 1261 -66 1264 -64
rect 1255 -76 1264 -66
rect 1222 -82 1229 -76
rect 1257 -82 1264 -76
rect 1266 -82 1271 -62
rect 1273 -69 1278 -62
rect 1316 -65 1321 -62
rect 1306 -68 1311 -65
rect 1273 -71 1280 -69
rect 1273 -73 1276 -71
rect 1278 -73 1280 -71
rect 1273 -75 1280 -73
rect 1284 -71 1291 -68
rect 1284 -73 1286 -71
rect 1288 -73 1291 -71
rect 1273 -82 1278 -75
rect 1284 -78 1291 -73
rect 1284 -80 1286 -78
rect 1288 -80 1291 -78
rect 1284 -82 1291 -80
rect 1293 -78 1301 -68
rect 1293 -80 1296 -78
rect 1298 -80 1301 -78
rect 1293 -82 1301 -80
rect 1303 -70 1311 -68
rect 1303 -72 1306 -70
rect 1308 -72 1311 -70
rect 1303 -75 1311 -72
rect 1313 -67 1321 -65
rect 1313 -69 1316 -67
rect 1318 -69 1321 -67
rect 1313 -75 1321 -69
rect 1323 -69 1328 -62
rect 1335 -65 1341 -63
rect 1335 -67 1337 -65
rect 1339 -67 1341 -65
rect 1335 -69 1341 -67
rect 1354 -65 1360 -63
rect 1401 -61 1408 -59
rect 1401 -63 1404 -61
rect 1406 -63 1408 -61
rect 1354 -67 1356 -65
rect 1358 -67 1360 -65
rect 1354 -69 1360 -67
rect 1323 -71 1330 -69
rect 1323 -73 1326 -71
rect 1328 -73 1330 -71
rect 1323 -75 1330 -73
rect 1303 -82 1308 -75
rect 1335 -76 1340 -69
rect 1356 -73 1360 -69
rect 1401 -69 1408 -63
rect 1383 -71 1390 -69
rect 1383 -73 1385 -71
rect 1387 -73 1390 -71
rect 1356 -76 1362 -73
rect 1335 -82 1342 -76
rect 1344 -78 1352 -76
rect 1344 -80 1347 -78
rect 1349 -80 1352 -78
rect 1344 -82 1352 -80
rect 1354 -82 1362 -76
rect 1364 -76 1369 -73
rect 1383 -75 1390 -73
rect 1364 -78 1371 -76
rect 1364 -80 1367 -78
rect 1369 -80 1371 -78
rect 1385 -80 1390 -75
rect 1392 -80 1397 -69
rect 1399 -71 1408 -69
rect 1425 -69 1430 -62
rect 1423 -71 1430 -69
rect 1399 -80 1410 -71
rect 1412 -73 1419 -71
rect 1412 -75 1415 -73
rect 1417 -75 1419 -73
rect 1423 -73 1425 -71
rect 1427 -73 1430 -71
rect 1423 -75 1430 -73
rect 1432 -65 1437 -62
rect 1432 -67 1440 -65
rect 1432 -69 1435 -67
rect 1437 -69 1440 -67
rect 1432 -75 1440 -69
rect 1442 -68 1447 -65
rect 1442 -70 1450 -68
rect 1442 -72 1445 -70
rect 1447 -72 1450 -70
rect 1442 -75 1450 -72
rect 1412 -77 1419 -75
rect 1412 -80 1417 -77
rect 1364 -82 1371 -80
rect 1445 -82 1450 -75
rect 1452 -78 1460 -68
rect 1452 -80 1455 -78
rect 1457 -80 1460 -78
rect 1452 -82 1460 -80
rect 1462 -71 1469 -68
rect 1475 -69 1480 -62
rect 1462 -73 1465 -71
rect 1467 -73 1469 -71
rect 1462 -78 1469 -73
rect 1473 -71 1480 -69
rect 1473 -73 1475 -71
rect 1477 -73 1480 -71
rect 1473 -75 1480 -73
rect 1462 -80 1465 -78
rect 1467 -80 1469 -78
rect 1462 -82 1469 -80
rect 1475 -82 1480 -75
rect 1482 -82 1487 -62
rect 1489 -64 1498 -62
rect 1489 -66 1492 -64
rect 1494 -66 1498 -64
rect 1489 -76 1498 -66
rect 1500 -69 1505 -62
rect 1515 -69 1520 -62
rect 1500 -71 1507 -69
rect 1500 -73 1503 -71
rect 1505 -73 1507 -71
rect 1500 -76 1507 -73
rect 1513 -71 1520 -69
rect 1513 -73 1515 -71
rect 1517 -73 1520 -71
rect 1513 -76 1520 -73
rect 1522 -64 1531 -62
rect 1522 -66 1526 -64
rect 1528 -66 1531 -64
rect 1522 -76 1531 -66
rect 1489 -82 1496 -76
rect 1524 -82 1531 -76
rect 1533 -82 1538 -62
rect 1540 -69 1545 -62
rect 1583 -65 1588 -62
rect 1573 -68 1578 -65
rect 1540 -71 1547 -69
rect 1540 -73 1543 -71
rect 1545 -73 1547 -71
rect 1540 -75 1547 -73
rect 1551 -71 1558 -68
rect 1551 -73 1553 -71
rect 1555 -73 1558 -71
rect 1540 -82 1545 -75
rect 1551 -78 1558 -73
rect 1551 -80 1553 -78
rect 1555 -80 1558 -78
rect 1551 -82 1558 -80
rect 1560 -78 1568 -68
rect 1560 -80 1563 -78
rect 1565 -80 1568 -78
rect 1560 -82 1568 -80
rect 1570 -70 1578 -68
rect 1570 -72 1573 -70
rect 1575 -72 1578 -70
rect 1570 -75 1578 -72
rect 1580 -67 1588 -65
rect 1580 -69 1583 -67
rect 1585 -69 1588 -67
rect 1580 -75 1588 -69
rect 1590 -69 1595 -62
rect 1602 -65 1608 -63
rect 1602 -67 1604 -65
rect 1606 -67 1608 -65
rect 1602 -69 1608 -67
rect 1621 -65 1627 -63
rect 1668 -61 1675 -59
rect 1668 -63 1671 -61
rect 1673 -63 1675 -61
rect 1621 -67 1623 -65
rect 1625 -67 1627 -65
rect 1621 -69 1627 -67
rect 1590 -71 1597 -69
rect 1590 -73 1593 -71
rect 1595 -73 1597 -71
rect 1590 -75 1597 -73
rect 1570 -82 1575 -75
rect 1602 -76 1607 -69
rect 1623 -73 1627 -69
rect 1668 -69 1675 -63
rect 1650 -71 1657 -69
rect 1650 -73 1652 -71
rect 1654 -73 1657 -71
rect 1623 -76 1629 -73
rect 1602 -82 1609 -76
rect 1611 -78 1619 -76
rect 1611 -80 1614 -78
rect 1616 -80 1619 -78
rect 1611 -82 1619 -80
rect 1621 -82 1629 -76
rect 1631 -76 1636 -73
rect 1650 -75 1657 -73
rect 1631 -78 1638 -76
rect 1631 -80 1634 -78
rect 1636 -80 1638 -78
rect 1652 -80 1657 -75
rect 1659 -80 1664 -69
rect 1666 -71 1675 -69
rect 1692 -69 1697 -62
rect 1690 -71 1697 -69
rect 1666 -80 1677 -71
rect 1679 -73 1686 -71
rect 1679 -75 1682 -73
rect 1684 -75 1686 -73
rect 1690 -73 1692 -71
rect 1694 -73 1697 -71
rect 1690 -75 1697 -73
rect 1699 -65 1704 -62
rect 1699 -67 1707 -65
rect 1699 -69 1702 -67
rect 1704 -69 1707 -67
rect 1699 -75 1707 -69
rect 1709 -68 1714 -65
rect 1709 -70 1717 -68
rect 1709 -72 1712 -70
rect 1714 -72 1717 -70
rect 1709 -75 1717 -72
rect 1679 -77 1686 -75
rect 1679 -80 1684 -77
rect 1631 -82 1638 -80
rect 1712 -82 1717 -75
rect 1719 -78 1727 -68
rect 1719 -80 1722 -78
rect 1724 -80 1727 -78
rect 1719 -82 1727 -80
rect 1729 -71 1736 -68
rect 1742 -69 1747 -62
rect 1729 -73 1732 -71
rect 1734 -73 1736 -71
rect 1729 -78 1736 -73
rect 1740 -71 1747 -69
rect 1740 -73 1742 -71
rect 1744 -73 1747 -71
rect 1740 -75 1747 -73
rect 1729 -80 1732 -78
rect 1734 -80 1736 -78
rect 1729 -82 1736 -80
rect 1742 -82 1747 -75
rect 1749 -82 1754 -62
rect 1756 -64 1765 -62
rect 1756 -66 1759 -64
rect 1761 -66 1765 -64
rect 1756 -76 1765 -66
rect 1767 -69 1772 -62
rect 1782 -69 1787 -62
rect 1767 -71 1774 -69
rect 1767 -73 1770 -71
rect 1772 -73 1774 -71
rect 1767 -76 1774 -73
rect 1780 -71 1787 -69
rect 1780 -73 1782 -71
rect 1784 -73 1787 -71
rect 1780 -76 1787 -73
rect 1789 -64 1798 -62
rect 1789 -66 1793 -64
rect 1795 -66 1798 -64
rect 1789 -76 1798 -66
rect 1756 -82 1763 -76
rect 1791 -82 1798 -76
rect 1800 -82 1805 -62
rect 1807 -69 1812 -62
rect 1850 -65 1855 -62
rect 1840 -68 1845 -65
rect 1807 -71 1814 -69
rect 1807 -73 1810 -71
rect 1812 -73 1814 -71
rect 1807 -75 1814 -73
rect 1818 -71 1825 -68
rect 1818 -73 1820 -71
rect 1822 -73 1825 -71
rect 1807 -82 1812 -75
rect 1818 -78 1825 -73
rect 1818 -80 1820 -78
rect 1822 -80 1825 -78
rect 1818 -82 1825 -80
rect 1827 -78 1835 -68
rect 1827 -80 1830 -78
rect 1832 -80 1835 -78
rect 1827 -82 1835 -80
rect 1837 -70 1845 -68
rect 1837 -72 1840 -70
rect 1842 -72 1845 -70
rect 1837 -75 1845 -72
rect 1847 -67 1855 -65
rect 1847 -69 1850 -67
rect 1852 -69 1855 -67
rect 1847 -75 1855 -69
rect 1857 -69 1862 -62
rect 1869 -65 1875 -63
rect 1869 -67 1871 -65
rect 1873 -67 1875 -65
rect 1869 -69 1875 -67
rect 1888 -65 1894 -63
rect 1888 -67 1890 -65
rect 1892 -67 1894 -65
rect 1888 -69 1894 -67
rect 1966 -61 1972 -59
rect 1966 -63 1968 -61
rect 1970 -63 1972 -61
rect 1966 -65 1972 -63
rect 1950 -68 1955 -65
rect 1857 -71 1864 -69
rect 1857 -73 1860 -71
rect 1862 -73 1864 -71
rect 1857 -75 1864 -73
rect 1837 -82 1842 -75
rect 1869 -76 1874 -69
rect 1890 -73 1894 -69
rect 1926 -70 1935 -68
rect 1926 -72 1928 -70
rect 1930 -72 1935 -70
rect 1926 -73 1935 -72
rect 1890 -76 1896 -73
rect 1869 -82 1876 -76
rect 1878 -78 1886 -76
rect 1878 -80 1881 -78
rect 1883 -80 1886 -78
rect 1878 -82 1886 -80
rect 1888 -82 1896 -76
rect 1898 -76 1903 -73
rect 1914 -76 1919 -73
rect 1898 -78 1905 -76
rect 1898 -80 1901 -78
rect 1903 -80 1905 -78
rect 1898 -82 1905 -80
rect 1912 -78 1919 -76
rect 1912 -80 1914 -78
rect 1916 -80 1919 -78
rect 1912 -82 1919 -80
rect 1921 -77 1935 -73
rect 1937 -73 1945 -68
rect 1937 -75 1940 -73
rect 1942 -75 1945 -73
rect 1937 -77 1945 -75
rect 1947 -71 1955 -68
rect 1947 -73 1950 -71
rect 1952 -73 1955 -71
rect 1947 -77 1955 -73
rect 1957 -77 1962 -65
rect 1964 -77 1972 -65
rect 1978 -69 1983 -62
rect 1976 -71 1983 -69
rect 1976 -73 1978 -71
rect 1980 -73 1983 -71
rect 1976 -75 1983 -73
rect 1985 -65 1990 -62
rect 1985 -67 1993 -65
rect 1985 -69 1988 -67
rect 1990 -69 1993 -67
rect 1985 -75 1993 -69
rect 1995 -68 2000 -65
rect 1995 -70 2003 -68
rect 1995 -72 1998 -70
rect 2000 -72 2003 -70
rect 1995 -75 2003 -72
rect 1921 -82 1926 -77
rect 1998 -82 2003 -75
rect 2005 -78 2013 -68
rect 2005 -80 2008 -78
rect 2010 -80 2013 -78
rect 2005 -82 2013 -80
rect 2015 -71 2022 -68
rect 2028 -69 2033 -62
rect 2015 -73 2018 -71
rect 2020 -73 2022 -71
rect 2015 -78 2022 -73
rect 2026 -71 2033 -69
rect 2026 -73 2028 -71
rect 2030 -73 2033 -71
rect 2026 -75 2033 -73
rect 2015 -80 2018 -78
rect 2020 -80 2022 -78
rect 2015 -82 2022 -80
rect 2028 -82 2033 -75
rect 2035 -82 2040 -62
rect 2042 -64 2051 -62
rect 2042 -66 2045 -64
rect 2047 -66 2051 -64
rect 2042 -76 2051 -66
rect 2053 -69 2058 -62
rect 2068 -69 2073 -62
rect 2053 -71 2060 -69
rect 2053 -73 2056 -71
rect 2058 -73 2060 -71
rect 2053 -76 2060 -73
rect 2066 -71 2073 -69
rect 2066 -73 2068 -71
rect 2070 -73 2073 -71
rect 2066 -76 2073 -73
rect 2075 -64 2084 -62
rect 2075 -66 2079 -64
rect 2081 -66 2084 -64
rect 2075 -76 2084 -66
rect 2042 -82 2049 -76
rect 2077 -82 2084 -76
rect 2086 -82 2091 -62
rect 2093 -69 2098 -62
rect 2136 -65 2141 -62
rect 2126 -68 2131 -65
rect 2093 -71 2100 -69
rect 2093 -73 2096 -71
rect 2098 -73 2100 -71
rect 2093 -75 2100 -73
rect 2104 -71 2111 -68
rect 2104 -73 2106 -71
rect 2108 -73 2111 -71
rect 2093 -82 2098 -75
rect 2104 -78 2111 -73
rect 2104 -80 2106 -78
rect 2108 -80 2111 -78
rect 2104 -82 2111 -80
rect 2113 -78 2121 -68
rect 2113 -80 2116 -78
rect 2118 -80 2121 -78
rect 2113 -82 2121 -80
rect 2123 -70 2131 -68
rect 2123 -72 2126 -70
rect 2128 -72 2131 -70
rect 2123 -75 2131 -72
rect 2133 -67 2141 -65
rect 2133 -69 2136 -67
rect 2138 -69 2141 -67
rect 2133 -75 2141 -69
rect 2143 -69 2148 -62
rect 2155 -65 2161 -63
rect 2155 -67 2157 -65
rect 2159 -67 2161 -65
rect 2155 -69 2161 -67
rect 2174 -65 2180 -63
rect 2174 -67 2176 -65
rect 2178 -67 2180 -65
rect 2174 -69 2180 -67
rect 2143 -71 2150 -69
rect 2143 -73 2146 -71
rect 2148 -73 2150 -71
rect 2143 -75 2150 -73
rect 2123 -82 2128 -75
rect 2155 -76 2160 -69
rect 2176 -73 2180 -69
rect 2210 -70 2216 -68
rect 2199 -72 2206 -70
rect 2176 -76 2182 -73
rect 2155 -82 2162 -76
rect 2164 -78 2172 -76
rect 2164 -80 2167 -78
rect 2169 -80 2172 -78
rect 2164 -82 2172 -80
rect 2174 -82 2182 -76
rect 2184 -76 2189 -73
rect 2199 -74 2201 -72
rect 2203 -74 2206 -72
rect 2199 -76 2206 -74
rect 2208 -72 2216 -70
rect 2208 -74 2211 -72
rect 2213 -74 2216 -72
rect 2208 -76 2216 -74
rect 2218 -76 2223 -68
rect 2225 -70 2233 -68
rect 2225 -72 2228 -70
rect 2230 -72 2233 -70
rect 2225 -76 2233 -72
rect 2235 -76 2240 -68
rect 2242 -70 2250 -68
rect 2242 -72 2245 -70
rect 2247 -72 2250 -70
rect 2242 -76 2250 -72
rect 2184 -78 2191 -76
rect 2184 -80 2187 -78
rect 2189 -80 2191 -78
rect 2184 -82 2191 -80
rect 2245 -77 2250 -76
rect 2252 -71 2257 -68
rect 2278 -70 2284 -68
rect 2252 -73 2259 -71
rect 2252 -75 2255 -73
rect 2257 -75 2259 -73
rect 2252 -77 2259 -75
rect 2267 -72 2274 -70
rect 2267 -74 2269 -72
rect 2271 -74 2274 -72
rect 2267 -76 2274 -74
rect 2276 -72 2284 -70
rect 2276 -74 2279 -72
rect 2281 -74 2284 -72
rect 2276 -76 2284 -74
rect 2286 -76 2291 -68
rect 2293 -70 2301 -68
rect 2293 -72 2296 -70
rect 2298 -72 2301 -70
rect 2293 -76 2301 -72
rect 2303 -76 2308 -68
rect 2310 -70 2318 -68
rect 2310 -72 2313 -70
rect 2315 -72 2318 -70
rect 2310 -76 2318 -72
rect 2313 -77 2318 -76
rect 2320 -71 2325 -68
rect 2320 -73 2327 -71
rect 2320 -75 2323 -73
rect 2325 -75 2327 -73
rect 2320 -77 2327 -75
rect 10 -181 15 -176
rect 8 -183 15 -181
rect 8 -185 10 -183
rect 12 -185 15 -183
rect 8 -187 15 -185
rect 17 -187 22 -176
rect 24 -185 35 -176
rect 37 -179 42 -176
rect 37 -181 44 -179
rect 50 -181 55 -176
rect 37 -183 40 -181
rect 42 -183 44 -181
rect 37 -185 44 -183
rect 48 -183 55 -181
rect 48 -185 50 -183
rect 52 -185 55 -183
rect 24 -187 33 -185
rect 26 -193 33 -187
rect 48 -187 55 -185
rect 57 -187 62 -176
rect 64 -185 75 -176
rect 77 -179 82 -176
rect 77 -181 84 -179
rect 110 -181 115 -174
rect 77 -183 80 -181
rect 82 -183 84 -181
rect 77 -185 84 -183
rect 88 -183 95 -181
rect 88 -185 90 -183
rect 92 -185 95 -183
rect 64 -187 73 -185
rect 26 -195 29 -193
rect 31 -195 33 -193
rect 26 -197 33 -195
rect 66 -193 73 -187
rect 88 -187 95 -185
rect 66 -195 69 -193
rect 71 -195 73 -193
rect 66 -197 73 -195
rect 90 -194 95 -187
rect 97 -187 105 -181
rect 97 -189 100 -187
rect 102 -189 105 -187
rect 97 -191 105 -189
rect 107 -184 115 -181
rect 107 -186 110 -184
rect 112 -186 115 -184
rect 107 -188 115 -186
rect 117 -176 125 -174
rect 117 -178 120 -176
rect 122 -178 125 -176
rect 117 -188 125 -178
rect 127 -176 134 -174
rect 127 -178 130 -176
rect 132 -178 134 -176
rect 127 -183 134 -178
rect 140 -181 145 -174
rect 127 -185 130 -183
rect 132 -185 134 -183
rect 127 -188 134 -185
rect 138 -183 145 -181
rect 138 -185 140 -183
rect 142 -185 145 -183
rect 138 -187 145 -185
rect 107 -191 112 -188
rect 97 -194 102 -191
rect 140 -194 145 -187
rect 147 -194 152 -174
rect 154 -180 161 -174
rect 189 -180 196 -174
rect 154 -190 163 -180
rect 154 -192 157 -190
rect 159 -192 163 -190
rect 154 -194 163 -192
rect 165 -183 172 -180
rect 165 -185 168 -183
rect 170 -185 172 -183
rect 165 -187 172 -185
rect 178 -183 185 -180
rect 178 -185 180 -183
rect 182 -185 185 -183
rect 178 -187 185 -185
rect 165 -194 170 -187
rect 180 -194 185 -187
rect 187 -190 196 -180
rect 187 -192 191 -190
rect 193 -192 196 -190
rect 187 -194 196 -192
rect 198 -194 203 -174
rect 205 -181 210 -174
rect 216 -176 223 -174
rect 216 -178 218 -176
rect 220 -178 223 -176
rect 205 -183 212 -181
rect 205 -185 208 -183
rect 210 -185 212 -183
rect 205 -187 212 -185
rect 216 -183 223 -178
rect 216 -185 218 -183
rect 220 -185 223 -183
rect 205 -194 210 -187
rect 216 -188 223 -185
rect 225 -176 233 -174
rect 225 -178 228 -176
rect 230 -178 233 -176
rect 225 -188 233 -178
rect 235 -181 240 -174
rect 267 -180 274 -174
rect 276 -176 284 -174
rect 276 -178 279 -176
rect 281 -178 284 -176
rect 276 -180 284 -178
rect 286 -180 294 -174
rect 235 -184 243 -181
rect 235 -186 238 -184
rect 240 -186 243 -184
rect 235 -188 243 -186
rect 238 -191 243 -188
rect 245 -187 253 -181
rect 245 -189 248 -187
rect 250 -189 253 -187
rect 245 -191 253 -189
rect 248 -194 253 -191
rect 255 -183 262 -181
rect 255 -185 258 -183
rect 260 -185 262 -183
rect 255 -187 262 -185
rect 267 -187 272 -180
rect 288 -183 294 -180
rect 296 -176 303 -174
rect 296 -178 299 -176
rect 301 -178 303 -176
rect 296 -180 303 -178
rect 296 -183 301 -180
rect 317 -181 322 -176
rect 315 -183 322 -181
rect 288 -187 292 -183
rect 255 -194 260 -187
rect 267 -189 273 -187
rect 267 -191 269 -189
rect 271 -191 273 -189
rect 267 -193 273 -191
rect 286 -189 292 -187
rect 315 -185 317 -183
rect 319 -185 322 -183
rect 315 -187 322 -185
rect 324 -187 329 -176
rect 331 -185 342 -176
rect 344 -179 349 -176
rect 344 -181 351 -179
rect 377 -181 382 -174
rect 344 -183 347 -181
rect 349 -183 351 -181
rect 344 -185 351 -183
rect 355 -183 362 -181
rect 355 -185 357 -183
rect 359 -185 362 -183
rect 331 -187 340 -185
rect 286 -191 288 -189
rect 290 -191 292 -189
rect 286 -193 292 -191
rect 333 -193 340 -187
rect 355 -187 362 -185
rect 333 -195 336 -193
rect 338 -195 340 -193
rect 333 -197 340 -195
rect 357 -194 362 -187
rect 364 -187 372 -181
rect 364 -189 367 -187
rect 369 -189 372 -187
rect 364 -191 372 -189
rect 374 -184 382 -181
rect 374 -186 377 -184
rect 379 -186 382 -184
rect 374 -188 382 -186
rect 384 -176 392 -174
rect 384 -178 387 -176
rect 389 -178 392 -176
rect 384 -188 392 -178
rect 394 -176 401 -174
rect 394 -178 397 -176
rect 399 -178 401 -176
rect 394 -183 401 -178
rect 407 -181 412 -174
rect 394 -185 397 -183
rect 399 -185 401 -183
rect 394 -188 401 -185
rect 405 -183 412 -181
rect 405 -185 407 -183
rect 409 -185 412 -183
rect 405 -187 412 -185
rect 374 -191 379 -188
rect 364 -194 369 -191
rect 407 -194 412 -187
rect 414 -194 419 -174
rect 421 -180 428 -174
rect 456 -180 463 -174
rect 421 -190 430 -180
rect 421 -192 424 -190
rect 426 -192 430 -190
rect 421 -194 430 -192
rect 432 -183 439 -180
rect 432 -185 435 -183
rect 437 -185 439 -183
rect 432 -187 439 -185
rect 445 -183 452 -180
rect 445 -185 447 -183
rect 449 -185 452 -183
rect 445 -187 452 -185
rect 432 -194 437 -187
rect 447 -194 452 -187
rect 454 -190 463 -180
rect 454 -192 458 -190
rect 460 -192 463 -190
rect 454 -194 463 -192
rect 465 -194 470 -174
rect 472 -181 477 -174
rect 483 -176 490 -174
rect 483 -178 485 -176
rect 487 -178 490 -176
rect 472 -183 479 -181
rect 472 -185 475 -183
rect 477 -185 479 -183
rect 472 -187 479 -185
rect 483 -183 490 -178
rect 483 -185 485 -183
rect 487 -185 490 -183
rect 472 -194 477 -187
rect 483 -188 490 -185
rect 492 -176 500 -174
rect 492 -178 495 -176
rect 497 -178 500 -176
rect 492 -188 500 -178
rect 502 -181 507 -174
rect 534 -180 541 -174
rect 543 -176 551 -174
rect 543 -178 546 -176
rect 548 -178 551 -176
rect 543 -180 551 -178
rect 553 -180 561 -174
rect 502 -184 510 -181
rect 502 -186 505 -184
rect 507 -186 510 -184
rect 502 -188 510 -186
rect 505 -191 510 -188
rect 512 -187 520 -181
rect 512 -189 515 -187
rect 517 -189 520 -187
rect 512 -191 520 -189
rect 515 -194 520 -191
rect 522 -183 529 -181
rect 522 -185 525 -183
rect 527 -185 529 -183
rect 522 -187 529 -185
rect 534 -187 539 -180
rect 555 -183 561 -180
rect 563 -176 570 -174
rect 563 -178 566 -176
rect 568 -178 570 -176
rect 563 -180 570 -178
rect 563 -183 568 -180
rect 584 -181 589 -176
rect 582 -183 589 -181
rect 555 -187 559 -183
rect 522 -194 527 -187
rect 534 -189 540 -187
rect 534 -191 536 -189
rect 538 -191 540 -189
rect 534 -193 540 -191
rect 553 -189 559 -187
rect 582 -185 584 -183
rect 586 -185 589 -183
rect 582 -187 589 -185
rect 591 -187 596 -176
rect 598 -185 609 -176
rect 611 -179 616 -176
rect 611 -181 618 -179
rect 644 -181 649 -174
rect 611 -183 614 -181
rect 616 -183 618 -181
rect 611 -185 618 -183
rect 622 -183 629 -181
rect 622 -185 624 -183
rect 626 -185 629 -183
rect 598 -187 607 -185
rect 553 -191 555 -189
rect 557 -191 559 -189
rect 553 -193 559 -191
rect 600 -193 607 -187
rect 622 -187 629 -185
rect 600 -195 603 -193
rect 605 -195 607 -193
rect 600 -197 607 -195
rect 624 -194 629 -187
rect 631 -187 639 -181
rect 631 -189 634 -187
rect 636 -189 639 -187
rect 631 -191 639 -189
rect 641 -184 649 -181
rect 641 -186 644 -184
rect 646 -186 649 -184
rect 641 -188 649 -186
rect 651 -176 659 -174
rect 651 -178 654 -176
rect 656 -178 659 -176
rect 651 -188 659 -178
rect 661 -176 668 -174
rect 661 -178 664 -176
rect 666 -178 668 -176
rect 661 -183 668 -178
rect 674 -181 679 -174
rect 661 -185 664 -183
rect 666 -185 668 -183
rect 661 -188 668 -185
rect 672 -183 679 -181
rect 672 -185 674 -183
rect 676 -185 679 -183
rect 672 -187 679 -185
rect 641 -191 646 -188
rect 631 -194 636 -191
rect 674 -194 679 -187
rect 681 -194 686 -174
rect 688 -180 695 -174
rect 723 -180 730 -174
rect 688 -190 697 -180
rect 688 -192 691 -190
rect 693 -192 697 -190
rect 688 -194 697 -192
rect 699 -183 706 -180
rect 699 -185 702 -183
rect 704 -185 706 -183
rect 699 -187 706 -185
rect 712 -183 719 -180
rect 712 -185 714 -183
rect 716 -185 719 -183
rect 712 -187 719 -185
rect 699 -194 704 -187
rect 714 -194 719 -187
rect 721 -190 730 -180
rect 721 -192 725 -190
rect 727 -192 730 -190
rect 721 -194 730 -192
rect 732 -194 737 -174
rect 739 -181 744 -174
rect 750 -176 757 -174
rect 750 -178 752 -176
rect 754 -178 757 -176
rect 739 -183 746 -181
rect 739 -185 742 -183
rect 744 -185 746 -183
rect 739 -187 746 -185
rect 750 -183 757 -178
rect 750 -185 752 -183
rect 754 -185 757 -183
rect 739 -194 744 -187
rect 750 -188 757 -185
rect 759 -176 767 -174
rect 759 -178 762 -176
rect 764 -178 767 -176
rect 759 -188 767 -178
rect 769 -181 774 -174
rect 801 -180 808 -174
rect 810 -176 818 -174
rect 810 -178 813 -176
rect 815 -178 818 -176
rect 810 -180 818 -178
rect 820 -180 828 -174
rect 769 -184 777 -181
rect 769 -186 772 -184
rect 774 -186 777 -184
rect 769 -188 777 -186
rect 772 -191 777 -188
rect 779 -187 787 -181
rect 779 -189 782 -187
rect 784 -189 787 -187
rect 779 -191 787 -189
rect 782 -194 787 -191
rect 789 -183 796 -181
rect 789 -185 792 -183
rect 794 -185 796 -183
rect 789 -187 796 -185
rect 801 -187 806 -180
rect 822 -183 828 -180
rect 830 -176 837 -174
rect 830 -178 833 -176
rect 835 -178 837 -176
rect 830 -180 837 -178
rect 830 -183 835 -180
rect 851 -181 856 -176
rect 849 -183 856 -181
rect 822 -187 826 -183
rect 789 -194 794 -187
rect 801 -189 807 -187
rect 801 -191 803 -189
rect 805 -191 807 -189
rect 801 -193 807 -191
rect 820 -189 826 -187
rect 849 -185 851 -183
rect 853 -185 856 -183
rect 849 -187 856 -185
rect 858 -187 863 -176
rect 865 -185 876 -176
rect 878 -179 883 -176
rect 878 -181 885 -179
rect 911 -181 916 -174
rect 878 -183 881 -181
rect 883 -183 885 -181
rect 878 -185 885 -183
rect 889 -183 896 -181
rect 889 -185 891 -183
rect 893 -185 896 -183
rect 865 -187 874 -185
rect 820 -191 822 -189
rect 824 -191 826 -189
rect 820 -193 826 -191
rect 867 -193 874 -187
rect 889 -187 896 -185
rect 867 -195 870 -193
rect 872 -195 874 -193
rect 867 -197 874 -195
rect 891 -194 896 -187
rect 898 -187 906 -181
rect 898 -189 901 -187
rect 903 -189 906 -187
rect 898 -191 906 -189
rect 908 -184 916 -181
rect 908 -186 911 -184
rect 913 -186 916 -184
rect 908 -188 916 -186
rect 918 -176 926 -174
rect 918 -178 921 -176
rect 923 -178 926 -176
rect 918 -188 926 -178
rect 928 -176 935 -174
rect 928 -178 931 -176
rect 933 -178 935 -176
rect 928 -183 935 -178
rect 941 -181 946 -174
rect 928 -185 931 -183
rect 933 -185 935 -183
rect 928 -188 935 -185
rect 939 -183 946 -181
rect 939 -185 941 -183
rect 943 -185 946 -183
rect 939 -187 946 -185
rect 908 -191 913 -188
rect 898 -194 903 -191
rect 941 -194 946 -187
rect 948 -194 953 -174
rect 955 -180 962 -174
rect 990 -180 997 -174
rect 955 -190 964 -180
rect 955 -192 958 -190
rect 960 -192 964 -190
rect 955 -194 964 -192
rect 966 -183 973 -180
rect 966 -185 969 -183
rect 971 -185 973 -183
rect 966 -187 973 -185
rect 979 -183 986 -180
rect 979 -185 981 -183
rect 983 -185 986 -183
rect 979 -187 986 -185
rect 966 -194 971 -187
rect 981 -194 986 -187
rect 988 -190 997 -180
rect 988 -192 992 -190
rect 994 -192 997 -190
rect 988 -194 997 -192
rect 999 -194 1004 -174
rect 1006 -181 1011 -174
rect 1017 -176 1024 -174
rect 1017 -178 1019 -176
rect 1021 -178 1024 -176
rect 1006 -183 1013 -181
rect 1006 -185 1009 -183
rect 1011 -185 1013 -183
rect 1006 -187 1013 -185
rect 1017 -183 1024 -178
rect 1017 -185 1019 -183
rect 1021 -185 1024 -183
rect 1006 -194 1011 -187
rect 1017 -188 1024 -185
rect 1026 -176 1034 -174
rect 1026 -178 1029 -176
rect 1031 -178 1034 -176
rect 1026 -188 1034 -178
rect 1036 -181 1041 -174
rect 1068 -180 1075 -174
rect 1077 -176 1085 -174
rect 1077 -178 1080 -176
rect 1082 -178 1085 -176
rect 1077 -180 1085 -178
rect 1087 -180 1095 -174
rect 1036 -184 1044 -181
rect 1036 -186 1039 -184
rect 1041 -186 1044 -184
rect 1036 -188 1044 -186
rect 1039 -191 1044 -188
rect 1046 -187 1054 -181
rect 1046 -189 1049 -187
rect 1051 -189 1054 -187
rect 1046 -191 1054 -189
rect 1049 -194 1054 -191
rect 1056 -183 1063 -181
rect 1056 -185 1059 -183
rect 1061 -185 1063 -183
rect 1056 -187 1063 -185
rect 1068 -187 1073 -180
rect 1089 -183 1095 -180
rect 1097 -176 1104 -174
rect 1097 -178 1100 -176
rect 1102 -178 1104 -176
rect 1097 -180 1104 -178
rect 1097 -183 1102 -180
rect 1118 -181 1123 -176
rect 1116 -183 1123 -181
rect 1089 -187 1093 -183
rect 1056 -194 1061 -187
rect 1068 -189 1074 -187
rect 1068 -191 1070 -189
rect 1072 -191 1074 -189
rect 1068 -193 1074 -191
rect 1087 -189 1093 -187
rect 1116 -185 1118 -183
rect 1120 -185 1123 -183
rect 1116 -187 1123 -185
rect 1125 -187 1130 -176
rect 1132 -185 1143 -176
rect 1145 -179 1150 -176
rect 1145 -181 1152 -179
rect 1178 -181 1183 -174
rect 1145 -183 1148 -181
rect 1150 -183 1152 -181
rect 1145 -185 1152 -183
rect 1156 -183 1163 -181
rect 1156 -185 1158 -183
rect 1160 -185 1163 -183
rect 1132 -187 1141 -185
rect 1087 -191 1089 -189
rect 1091 -191 1093 -189
rect 1087 -193 1093 -191
rect 1134 -193 1141 -187
rect 1156 -187 1163 -185
rect 1134 -195 1137 -193
rect 1139 -195 1141 -193
rect 1134 -197 1141 -195
rect 1158 -194 1163 -187
rect 1165 -187 1173 -181
rect 1165 -189 1168 -187
rect 1170 -189 1173 -187
rect 1165 -191 1173 -189
rect 1175 -184 1183 -181
rect 1175 -186 1178 -184
rect 1180 -186 1183 -184
rect 1175 -188 1183 -186
rect 1185 -176 1193 -174
rect 1185 -178 1188 -176
rect 1190 -178 1193 -176
rect 1185 -188 1193 -178
rect 1195 -176 1202 -174
rect 1195 -178 1198 -176
rect 1200 -178 1202 -176
rect 1195 -183 1202 -178
rect 1208 -181 1213 -174
rect 1195 -185 1198 -183
rect 1200 -185 1202 -183
rect 1195 -188 1202 -185
rect 1206 -183 1213 -181
rect 1206 -185 1208 -183
rect 1210 -185 1213 -183
rect 1206 -187 1213 -185
rect 1175 -191 1180 -188
rect 1165 -194 1170 -191
rect 1208 -194 1213 -187
rect 1215 -194 1220 -174
rect 1222 -180 1229 -174
rect 1257 -180 1264 -174
rect 1222 -190 1231 -180
rect 1222 -192 1225 -190
rect 1227 -192 1231 -190
rect 1222 -194 1231 -192
rect 1233 -183 1240 -180
rect 1233 -185 1236 -183
rect 1238 -185 1240 -183
rect 1233 -187 1240 -185
rect 1246 -183 1253 -180
rect 1246 -185 1248 -183
rect 1250 -185 1253 -183
rect 1246 -187 1253 -185
rect 1233 -194 1238 -187
rect 1248 -194 1253 -187
rect 1255 -190 1264 -180
rect 1255 -192 1259 -190
rect 1261 -192 1264 -190
rect 1255 -194 1264 -192
rect 1266 -194 1271 -174
rect 1273 -181 1278 -174
rect 1284 -176 1291 -174
rect 1284 -178 1286 -176
rect 1288 -178 1291 -176
rect 1273 -183 1280 -181
rect 1273 -185 1276 -183
rect 1278 -185 1280 -183
rect 1273 -187 1280 -185
rect 1284 -183 1291 -178
rect 1284 -185 1286 -183
rect 1288 -185 1291 -183
rect 1273 -194 1278 -187
rect 1284 -188 1291 -185
rect 1293 -176 1301 -174
rect 1293 -178 1296 -176
rect 1298 -178 1301 -176
rect 1293 -188 1301 -178
rect 1303 -181 1308 -174
rect 1335 -180 1342 -174
rect 1344 -176 1352 -174
rect 1344 -178 1347 -176
rect 1349 -178 1352 -176
rect 1344 -180 1352 -178
rect 1354 -180 1362 -174
rect 1303 -184 1311 -181
rect 1303 -186 1306 -184
rect 1308 -186 1311 -184
rect 1303 -188 1311 -186
rect 1306 -191 1311 -188
rect 1313 -187 1321 -181
rect 1313 -189 1316 -187
rect 1318 -189 1321 -187
rect 1313 -191 1321 -189
rect 1316 -194 1321 -191
rect 1323 -183 1330 -181
rect 1323 -185 1326 -183
rect 1328 -185 1330 -183
rect 1323 -187 1330 -185
rect 1335 -187 1340 -180
rect 1356 -183 1362 -180
rect 1364 -176 1371 -174
rect 1364 -178 1367 -176
rect 1369 -178 1371 -176
rect 1364 -180 1371 -178
rect 1364 -183 1369 -180
rect 1385 -181 1390 -176
rect 1383 -183 1390 -181
rect 1356 -187 1360 -183
rect 1323 -194 1328 -187
rect 1335 -189 1341 -187
rect 1335 -191 1337 -189
rect 1339 -191 1341 -189
rect 1335 -193 1341 -191
rect 1354 -189 1360 -187
rect 1383 -185 1385 -183
rect 1387 -185 1390 -183
rect 1383 -187 1390 -185
rect 1392 -187 1397 -176
rect 1399 -185 1410 -176
rect 1412 -179 1417 -176
rect 1412 -181 1419 -179
rect 1445 -181 1450 -174
rect 1412 -183 1415 -181
rect 1417 -183 1419 -181
rect 1412 -185 1419 -183
rect 1423 -183 1430 -181
rect 1423 -185 1425 -183
rect 1427 -185 1430 -183
rect 1399 -187 1408 -185
rect 1354 -191 1356 -189
rect 1358 -191 1360 -189
rect 1354 -193 1360 -191
rect 1401 -193 1408 -187
rect 1423 -187 1430 -185
rect 1401 -195 1404 -193
rect 1406 -195 1408 -193
rect 1401 -197 1408 -195
rect 1425 -194 1430 -187
rect 1432 -187 1440 -181
rect 1432 -189 1435 -187
rect 1437 -189 1440 -187
rect 1432 -191 1440 -189
rect 1442 -184 1450 -181
rect 1442 -186 1445 -184
rect 1447 -186 1450 -184
rect 1442 -188 1450 -186
rect 1452 -176 1460 -174
rect 1452 -178 1455 -176
rect 1457 -178 1460 -176
rect 1452 -188 1460 -178
rect 1462 -176 1469 -174
rect 1462 -178 1465 -176
rect 1467 -178 1469 -176
rect 1462 -183 1469 -178
rect 1475 -181 1480 -174
rect 1462 -185 1465 -183
rect 1467 -185 1469 -183
rect 1462 -188 1469 -185
rect 1473 -183 1480 -181
rect 1473 -185 1475 -183
rect 1477 -185 1480 -183
rect 1473 -187 1480 -185
rect 1442 -191 1447 -188
rect 1432 -194 1437 -191
rect 1475 -194 1480 -187
rect 1482 -194 1487 -174
rect 1489 -180 1496 -174
rect 1524 -180 1531 -174
rect 1489 -190 1498 -180
rect 1489 -192 1492 -190
rect 1494 -192 1498 -190
rect 1489 -194 1498 -192
rect 1500 -183 1507 -180
rect 1500 -185 1503 -183
rect 1505 -185 1507 -183
rect 1500 -187 1507 -185
rect 1513 -183 1520 -180
rect 1513 -185 1515 -183
rect 1517 -185 1520 -183
rect 1513 -187 1520 -185
rect 1500 -194 1505 -187
rect 1515 -194 1520 -187
rect 1522 -190 1531 -180
rect 1522 -192 1526 -190
rect 1528 -192 1531 -190
rect 1522 -194 1531 -192
rect 1533 -194 1538 -174
rect 1540 -181 1545 -174
rect 1551 -176 1558 -174
rect 1551 -178 1553 -176
rect 1555 -178 1558 -176
rect 1540 -183 1547 -181
rect 1540 -185 1543 -183
rect 1545 -185 1547 -183
rect 1540 -187 1547 -185
rect 1551 -183 1558 -178
rect 1551 -185 1553 -183
rect 1555 -185 1558 -183
rect 1540 -194 1545 -187
rect 1551 -188 1558 -185
rect 1560 -176 1568 -174
rect 1560 -178 1563 -176
rect 1565 -178 1568 -176
rect 1560 -188 1568 -178
rect 1570 -181 1575 -174
rect 1602 -180 1609 -174
rect 1611 -176 1619 -174
rect 1611 -178 1614 -176
rect 1616 -178 1619 -176
rect 1611 -180 1619 -178
rect 1621 -180 1629 -174
rect 1570 -184 1578 -181
rect 1570 -186 1573 -184
rect 1575 -186 1578 -184
rect 1570 -188 1578 -186
rect 1573 -191 1578 -188
rect 1580 -187 1588 -181
rect 1580 -189 1583 -187
rect 1585 -189 1588 -187
rect 1580 -191 1588 -189
rect 1583 -194 1588 -191
rect 1590 -183 1597 -181
rect 1590 -185 1593 -183
rect 1595 -185 1597 -183
rect 1590 -187 1597 -185
rect 1602 -187 1607 -180
rect 1623 -183 1629 -180
rect 1631 -176 1638 -174
rect 1631 -178 1634 -176
rect 1636 -178 1638 -176
rect 1631 -180 1638 -178
rect 1631 -183 1636 -180
rect 1652 -181 1657 -176
rect 1650 -183 1657 -181
rect 1623 -187 1627 -183
rect 1590 -194 1595 -187
rect 1602 -189 1608 -187
rect 1602 -191 1604 -189
rect 1606 -191 1608 -189
rect 1602 -193 1608 -191
rect 1621 -189 1627 -187
rect 1650 -185 1652 -183
rect 1654 -185 1657 -183
rect 1650 -187 1657 -185
rect 1659 -187 1664 -176
rect 1666 -185 1677 -176
rect 1679 -179 1684 -176
rect 1679 -181 1686 -179
rect 1712 -181 1717 -174
rect 1679 -183 1682 -181
rect 1684 -183 1686 -181
rect 1679 -185 1686 -183
rect 1690 -183 1697 -181
rect 1690 -185 1692 -183
rect 1694 -185 1697 -183
rect 1666 -187 1675 -185
rect 1621 -191 1623 -189
rect 1625 -191 1627 -189
rect 1621 -193 1627 -191
rect 1668 -193 1675 -187
rect 1690 -187 1697 -185
rect 1668 -195 1671 -193
rect 1673 -195 1675 -193
rect 1668 -197 1675 -195
rect 1692 -194 1697 -187
rect 1699 -187 1707 -181
rect 1699 -189 1702 -187
rect 1704 -189 1707 -187
rect 1699 -191 1707 -189
rect 1709 -184 1717 -181
rect 1709 -186 1712 -184
rect 1714 -186 1717 -184
rect 1709 -188 1717 -186
rect 1719 -176 1727 -174
rect 1719 -178 1722 -176
rect 1724 -178 1727 -176
rect 1719 -188 1727 -178
rect 1729 -176 1736 -174
rect 1729 -178 1732 -176
rect 1734 -178 1736 -176
rect 1729 -183 1736 -178
rect 1742 -181 1747 -174
rect 1729 -185 1732 -183
rect 1734 -185 1736 -183
rect 1729 -188 1736 -185
rect 1740 -183 1747 -181
rect 1740 -185 1742 -183
rect 1744 -185 1747 -183
rect 1740 -187 1747 -185
rect 1709 -191 1714 -188
rect 1699 -194 1704 -191
rect 1742 -194 1747 -187
rect 1749 -194 1754 -174
rect 1756 -180 1763 -174
rect 1791 -180 1798 -174
rect 1756 -190 1765 -180
rect 1756 -192 1759 -190
rect 1761 -192 1765 -190
rect 1756 -194 1765 -192
rect 1767 -183 1774 -180
rect 1767 -185 1770 -183
rect 1772 -185 1774 -183
rect 1767 -187 1774 -185
rect 1780 -183 1787 -180
rect 1780 -185 1782 -183
rect 1784 -185 1787 -183
rect 1780 -187 1787 -185
rect 1767 -194 1772 -187
rect 1782 -194 1787 -187
rect 1789 -190 1798 -180
rect 1789 -192 1793 -190
rect 1795 -192 1798 -190
rect 1789 -194 1798 -192
rect 1800 -194 1805 -174
rect 1807 -181 1812 -174
rect 1818 -176 1825 -174
rect 1818 -178 1820 -176
rect 1822 -178 1825 -176
rect 1807 -183 1814 -181
rect 1807 -185 1810 -183
rect 1812 -185 1814 -183
rect 1807 -187 1814 -185
rect 1818 -183 1825 -178
rect 1818 -185 1820 -183
rect 1822 -185 1825 -183
rect 1807 -194 1812 -187
rect 1818 -188 1825 -185
rect 1827 -176 1835 -174
rect 1827 -178 1830 -176
rect 1832 -178 1835 -176
rect 1827 -188 1835 -178
rect 1837 -181 1842 -174
rect 1869 -180 1876 -174
rect 1878 -176 1886 -174
rect 1878 -178 1881 -176
rect 1883 -178 1886 -176
rect 1878 -180 1886 -178
rect 1888 -180 1896 -174
rect 1837 -184 1845 -181
rect 1837 -186 1840 -184
rect 1842 -186 1845 -184
rect 1837 -188 1845 -186
rect 1840 -191 1845 -188
rect 1847 -187 1855 -181
rect 1847 -189 1850 -187
rect 1852 -189 1855 -187
rect 1847 -191 1855 -189
rect 1850 -194 1855 -191
rect 1857 -183 1864 -181
rect 1857 -185 1860 -183
rect 1862 -185 1864 -183
rect 1857 -187 1864 -185
rect 1869 -187 1874 -180
rect 1890 -183 1896 -180
rect 1898 -176 1905 -174
rect 1898 -178 1901 -176
rect 1903 -178 1905 -176
rect 1898 -180 1905 -178
rect 1912 -176 1919 -174
rect 1912 -178 1914 -176
rect 1916 -178 1919 -176
rect 1912 -180 1919 -178
rect 1898 -183 1903 -180
rect 1914 -183 1919 -180
rect 1921 -179 1926 -174
rect 1921 -183 1935 -179
rect 1890 -187 1894 -183
rect 1857 -194 1862 -187
rect 1869 -189 1875 -187
rect 1869 -191 1871 -189
rect 1873 -191 1875 -189
rect 1869 -193 1875 -191
rect 1888 -189 1894 -187
rect 1926 -184 1935 -183
rect 1926 -186 1928 -184
rect 1930 -186 1935 -184
rect 1926 -188 1935 -186
rect 1937 -181 1945 -179
rect 1937 -183 1940 -181
rect 1942 -183 1945 -181
rect 1937 -188 1945 -183
rect 1947 -183 1955 -179
rect 1947 -185 1950 -183
rect 1952 -185 1955 -183
rect 1947 -188 1955 -185
rect 1888 -191 1890 -189
rect 1892 -191 1894 -189
rect 1888 -193 1894 -191
rect 1950 -191 1955 -188
rect 1957 -191 1962 -179
rect 1964 -191 1972 -179
rect 1998 -181 2003 -174
rect 1976 -183 1983 -181
rect 1976 -185 1978 -183
rect 1980 -185 1983 -183
rect 1976 -187 1983 -185
rect 1966 -193 1972 -191
rect 1966 -195 1968 -193
rect 1970 -195 1972 -193
rect 1978 -194 1983 -187
rect 1985 -187 1993 -181
rect 1985 -189 1988 -187
rect 1990 -189 1993 -187
rect 1985 -191 1993 -189
rect 1995 -184 2003 -181
rect 1995 -186 1998 -184
rect 2000 -186 2003 -184
rect 1995 -188 2003 -186
rect 2005 -176 2013 -174
rect 2005 -178 2008 -176
rect 2010 -178 2013 -176
rect 2005 -188 2013 -178
rect 2015 -176 2022 -174
rect 2015 -178 2018 -176
rect 2020 -178 2022 -176
rect 2015 -183 2022 -178
rect 2028 -181 2033 -174
rect 2015 -185 2018 -183
rect 2020 -185 2022 -183
rect 2015 -188 2022 -185
rect 2026 -183 2033 -181
rect 2026 -185 2028 -183
rect 2030 -185 2033 -183
rect 2026 -187 2033 -185
rect 1995 -191 2000 -188
rect 1985 -194 1990 -191
rect 1966 -197 1972 -195
rect 2028 -194 2033 -187
rect 2035 -194 2040 -174
rect 2042 -180 2049 -174
rect 2077 -180 2084 -174
rect 2042 -190 2051 -180
rect 2042 -192 2045 -190
rect 2047 -192 2051 -190
rect 2042 -194 2051 -192
rect 2053 -183 2060 -180
rect 2053 -185 2056 -183
rect 2058 -185 2060 -183
rect 2053 -187 2060 -185
rect 2066 -183 2073 -180
rect 2066 -185 2068 -183
rect 2070 -185 2073 -183
rect 2066 -187 2073 -185
rect 2053 -194 2058 -187
rect 2068 -194 2073 -187
rect 2075 -190 2084 -180
rect 2075 -192 2079 -190
rect 2081 -192 2084 -190
rect 2075 -194 2084 -192
rect 2086 -194 2091 -174
rect 2093 -181 2098 -174
rect 2104 -176 2111 -174
rect 2104 -178 2106 -176
rect 2108 -178 2111 -176
rect 2093 -183 2100 -181
rect 2093 -185 2096 -183
rect 2098 -185 2100 -183
rect 2093 -187 2100 -185
rect 2104 -183 2111 -178
rect 2104 -185 2106 -183
rect 2108 -185 2111 -183
rect 2093 -194 2098 -187
rect 2104 -188 2111 -185
rect 2113 -176 2121 -174
rect 2113 -178 2116 -176
rect 2118 -178 2121 -176
rect 2113 -188 2121 -178
rect 2123 -181 2128 -174
rect 2155 -180 2162 -174
rect 2164 -176 2172 -174
rect 2164 -178 2167 -176
rect 2169 -178 2172 -176
rect 2164 -180 2172 -178
rect 2174 -180 2182 -174
rect 2123 -184 2131 -181
rect 2123 -186 2126 -184
rect 2128 -186 2131 -184
rect 2123 -188 2131 -186
rect 2126 -191 2131 -188
rect 2133 -187 2141 -181
rect 2133 -189 2136 -187
rect 2138 -189 2141 -187
rect 2133 -191 2141 -189
rect 2136 -194 2141 -191
rect 2143 -183 2150 -181
rect 2143 -185 2146 -183
rect 2148 -185 2150 -183
rect 2143 -187 2150 -185
rect 2155 -187 2160 -180
rect 2176 -183 2182 -180
rect 2184 -176 2191 -174
rect 2184 -178 2187 -176
rect 2189 -178 2191 -176
rect 2184 -180 2191 -178
rect 2245 -180 2250 -179
rect 2184 -183 2189 -180
rect 2199 -182 2206 -180
rect 2176 -187 2180 -183
rect 2143 -194 2148 -187
rect 2155 -189 2161 -187
rect 2155 -191 2157 -189
rect 2159 -191 2161 -189
rect 2155 -193 2161 -191
rect 2174 -189 2180 -187
rect 2199 -184 2201 -182
rect 2203 -184 2206 -182
rect 2199 -186 2206 -184
rect 2208 -182 2216 -180
rect 2208 -184 2211 -182
rect 2213 -184 2216 -182
rect 2208 -186 2216 -184
rect 2174 -191 2176 -189
rect 2178 -191 2180 -189
rect 2174 -193 2180 -191
rect 2210 -188 2216 -186
rect 2218 -188 2223 -180
rect 2225 -184 2233 -180
rect 2225 -186 2228 -184
rect 2230 -186 2233 -184
rect 2225 -188 2233 -186
rect 2235 -188 2240 -180
rect 2242 -184 2250 -180
rect 2242 -186 2245 -184
rect 2247 -186 2250 -184
rect 2242 -188 2250 -186
rect 2252 -181 2259 -179
rect 2313 -180 2318 -179
rect 2252 -183 2255 -181
rect 2257 -183 2259 -181
rect 2252 -185 2259 -183
rect 2267 -182 2274 -180
rect 2267 -184 2269 -182
rect 2271 -184 2274 -182
rect 2252 -188 2257 -185
rect 2267 -186 2274 -184
rect 2276 -182 2284 -180
rect 2276 -184 2279 -182
rect 2281 -184 2284 -182
rect 2276 -186 2284 -184
rect 2278 -188 2284 -186
rect 2286 -188 2291 -180
rect 2293 -184 2301 -180
rect 2293 -186 2296 -184
rect 2298 -186 2301 -184
rect 2293 -188 2301 -186
rect 2303 -188 2308 -180
rect 2310 -184 2318 -180
rect 2310 -186 2313 -184
rect 2315 -186 2318 -184
rect 2310 -188 2318 -186
rect 2320 -181 2327 -179
rect 2320 -183 2323 -181
rect 2325 -183 2327 -181
rect 2320 -185 2327 -183
rect 2320 -188 2325 -185
rect 26 -205 33 -203
rect 26 -207 29 -205
rect 31 -207 33 -205
rect 26 -213 33 -207
rect 66 -205 73 -203
rect 66 -207 69 -205
rect 71 -207 73 -205
rect 8 -215 15 -213
rect 8 -217 10 -215
rect 12 -217 15 -215
rect 8 -219 15 -217
rect 10 -224 15 -219
rect 17 -224 22 -213
rect 24 -215 33 -213
rect 66 -213 73 -207
rect 48 -215 55 -213
rect 24 -224 35 -215
rect 37 -217 44 -215
rect 37 -219 40 -217
rect 42 -219 44 -217
rect 48 -217 50 -215
rect 52 -217 55 -215
rect 48 -219 55 -217
rect 37 -221 44 -219
rect 37 -224 42 -221
rect 50 -224 55 -219
rect 57 -224 62 -213
rect 64 -215 73 -213
rect 90 -213 95 -206
rect 88 -215 95 -213
rect 64 -224 75 -215
rect 77 -217 84 -215
rect 77 -219 80 -217
rect 82 -219 84 -217
rect 88 -217 90 -215
rect 92 -217 95 -215
rect 88 -219 95 -217
rect 97 -209 102 -206
rect 97 -211 105 -209
rect 97 -213 100 -211
rect 102 -213 105 -211
rect 97 -219 105 -213
rect 107 -212 112 -209
rect 107 -214 115 -212
rect 107 -216 110 -214
rect 112 -216 115 -214
rect 107 -219 115 -216
rect 77 -221 84 -219
rect 77 -224 82 -221
rect 110 -226 115 -219
rect 117 -222 125 -212
rect 117 -224 120 -222
rect 122 -224 125 -222
rect 117 -226 125 -224
rect 127 -215 134 -212
rect 140 -213 145 -206
rect 127 -217 130 -215
rect 132 -217 134 -215
rect 127 -222 134 -217
rect 138 -215 145 -213
rect 138 -217 140 -215
rect 142 -217 145 -215
rect 138 -219 145 -217
rect 127 -224 130 -222
rect 132 -224 134 -222
rect 127 -226 134 -224
rect 140 -226 145 -219
rect 147 -226 152 -206
rect 154 -208 163 -206
rect 154 -210 157 -208
rect 159 -210 163 -208
rect 154 -220 163 -210
rect 165 -213 170 -206
rect 180 -213 185 -206
rect 165 -215 172 -213
rect 165 -217 168 -215
rect 170 -217 172 -215
rect 165 -220 172 -217
rect 178 -215 185 -213
rect 178 -217 180 -215
rect 182 -217 185 -215
rect 178 -220 185 -217
rect 187 -208 196 -206
rect 187 -210 191 -208
rect 193 -210 196 -208
rect 187 -220 196 -210
rect 154 -226 161 -220
rect 189 -226 196 -220
rect 198 -226 203 -206
rect 205 -213 210 -206
rect 248 -209 253 -206
rect 238 -212 243 -209
rect 205 -215 212 -213
rect 205 -217 208 -215
rect 210 -217 212 -215
rect 205 -219 212 -217
rect 216 -215 223 -212
rect 216 -217 218 -215
rect 220 -217 223 -215
rect 205 -226 210 -219
rect 216 -222 223 -217
rect 216 -224 218 -222
rect 220 -224 223 -222
rect 216 -226 223 -224
rect 225 -222 233 -212
rect 225 -224 228 -222
rect 230 -224 233 -222
rect 225 -226 233 -224
rect 235 -214 243 -212
rect 235 -216 238 -214
rect 240 -216 243 -214
rect 235 -219 243 -216
rect 245 -211 253 -209
rect 245 -213 248 -211
rect 250 -213 253 -211
rect 245 -219 253 -213
rect 255 -213 260 -206
rect 267 -209 273 -207
rect 267 -211 269 -209
rect 271 -211 273 -209
rect 267 -213 273 -211
rect 286 -209 292 -207
rect 333 -205 340 -203
rect 333 -207 336 -205
rect 338 -207 340 -205
rect 286 -211 288 -209
rect 290 -211 292 -209
rect 286 -213 292 -211
rect 255 -215 262 -213
rect 255 -217 258 -215
rect 260 -217 262 -215
rect 255 -219 262 -217
rect 235 -226 240 -219
rect 267 -220 272 -213
rect 288 -217 292 -213
rect 333 -213 340 -207
rect 315 -215 322 -213
rect 315 -217 317 -215
rect 319 -217 322 -215
rect 288 -220 294 -217
rect 267 -226 274 -220
rect 276 -222 284 -220
rect 276 -224 279 -222
rect 281 -224 284 -222
rect 276 -226 284 -224
rect 286 -226 294 -220
rect 296 -220 301 -217
rect 315 -219 322 -217
rect 296 -222 303 -220
rect 296 -224 299 -222
rect 301 -224 303 -222
rect 317 -224 322 -219
rect 324 -224 329 -213
rect 331 -215 340 -213
rect 357 -213 362 -206
rect 355 -215 362 -213
rect 331 -224 342 -215
rect 344 -217 351 -215
rect 344 -219 347 -217
rect 349 -219 351 -217
rect 355 -217 357 -215
rect 359 -217 362 -215
rect 355 -219 362 -217
rect 364 -209 369 -206
rect 364 -211 372 -209
rect 364 -213 367 -211
rect 369 -213 372 -211
rect 364 -219 372 -213
rect 374 -212 379 -209
rect 374 -214 382 -212
rect 374 -216 377 -214
rect 379 -216 382 -214
rect 374 -219 382 -216
rect 344 -221 351 -219
rect 344 -224 349 -221
rect 296 -226 303 -224
rect 377 -226 382 -219
rect 384 -222 392 -212
rect 384 -224 387 -222
rect 389 -224 392 -222
rect 384 -226 392 -224
rect 394 -215 401 -212
rect 407 -213 412 -206
rect 394 -217 397 -215
rect 399 -217 401 -215
rect 394 -222 401 -217
rect 405 -215 412 -213
rect 405 -217 407 -215
rect 409 -217 412 -215
rect 405 -219 412 -217
rect 394 -224 397 -222
rect 399 -224 401 -222
rect 394 -226 401 -224
rect 407 -226 412 -219
rect 414 -226 419 -206
rect 421 -208 430 -206
rect 421 -210 424 -208
rect 426 -210 430 -208
rect 421 -220 430 -210
rect 432 -213 437 -206
rect 447 -213 452 -206
rect 432 -215 439 -213
rect 432 -217 435 -215
rect 437 -217 439 -215
rect 432 -220 439 -217
rect 445 -215 452 -213
rect 445 -217 447 -215
rect 449 -217 452 -215
rect 445 -220 452 -217
rect 454 -208 463 -206
rect 454 -210 458 -208
rect 460 -210 463 -208
rect 454 -220 463 -210
rect 421 -226 428 -220
rect 456 -226 463 -220
rect 465 -226 470 -206
rect 472 -213 477 -206
rect 515 -209 520 -206
rect 505 -212 510 -209
rect 472 -215 479 -213
rect 472 -217 475 -215
rect 477 -217 479 -215
rect 472 -219 479 -217
rect 483 -215 490 -212
rect 483 -217 485 -215
rect 487 -217 490 -215
rect 472 -226 477 -219
rect 483 -222 490 -217
rect 483 -224 485 -222
rect 487 -224 490 -222
rect 483 -226 490 -224
rect 492 -222 500 -212
rect 492 -224 495 -222
rect 497 -224 500 -222
rect 492 -226 500 -224
rect 502 -214 510 -212
rect 502 -216 505 -214
rect 507 -216 510 -214
rect 502 -219 510 -216
rect 512 -211 520 -209
rect 512 -213 515 -211
rect 517 -213 520 -211
rect 512 -219 520 -213
rect 522 -213 527 -206
rect 534 -209 540 -207
rect 534 -211 536 -209
rect 538 -211 540 -209
rect 534 -213 540 -211
rect 553 -209 559 -207
rect 600 -205 607 -203
rect 600 -207 603 -205
rect 605 -207 607 -205
rect 553 -211 555 -209
rect 557 -211 559 -209
rect 553 -213 559 -211
rect 522 -215 529 -213
rect 522 -217 525 -215
rect 527 -217 529 -215
rect 522 -219 529 -217
rect 502 -226 507 -219
rect 534 -220 539 -213
rect 555 -217 559 -213
rect 600 -213 607 -207
rect 582 -215 589 -213
rect 582 -217 584 -215
rect 586 -217 589 -215
rect 555 -220 561 -217
rect 534 -226 541 -220
rect 543 -222 551 -220
rect 543 -224 546 -222
rect 548 -224 551 -222
rect 543 -226 551 -224
rect 553 -226 561 -220
rect 563 -220 568 -217
rect 582 -219 589 -217
rect 563 -222 570 -220
rect 563 -224 566 -222
rect 568 -224 570 -222
rect 584 -224 589 -219
rect 591 -224 596 -213
rect 598 -215 607 -213
rect 624 -213 629 -206
rect 622 -215 629 -213
rect 598 -224 609 -215
rect 611 -217 618 -215
rect 611 -219 614 -217
rect 616 -219 618 -217
rect 622 -217 624 -215
rect 626 -217 629 -215
rect 622 -219 629 -217
rect 631 -209 636 -206
rect 631 -211 639 -209
rect 631 -213 634 -211
rect 636 -213 639 -211
rect 631 -219 639 -213
rect 641 -212 646 -209
rect 641 -214 649 -212
rect 641 -216 644 -214
rect 646 -216 649 -214
rect 641 -219 649 -216
rect 611 -221 618 -219
rect 611 -224 616 -221
rect 563 -226 570 -224
rect 644 -226 649 -219
rect 651 -222 659 -212
rect 651 -224 654 -222
rect 656 -224 659 -222
rect 651 -226 659 -224
rect 661 -215 668 -212
rect 674 -213 679 -206
rect 661 -217 664 -215
rect 666 -217 668 -215
rect 661 -222 668 -217
rect 672 -215 679 -213
rect 672 -217 674 -215
rect 676 -217 679 -215
rect 672 -219 679 -217
rect 661 -224 664 -222
rect 666 -224 668 -222
rect 661 -226 668 -224
rect 674 -226 679 -219
rect 681 -226 686 -206
rect 688 -208 697 -206
rect 688 -210 691 -208
rect 693 -210 697 -208
rect 688 -220 697 -210
rect 699 -213 704 -206
rect 714 -213 719 -206
rect 699 -215 706 -213
rect 699 -217 702 -215
rect 704 -217 706 -215
rect 699 -220 706 -217
rect 712 -215 719 -213
rect 712 -217 714 -215
rect 716 -217 719 -215
rect 712 -220 719 -217
rect 721 -208 730 -206
rect 721 -210 725 -208
rect 727 -210 730 -208
rect 721 -220 730 -210
rect 688 -226 695 -220
rect 723 -226 730 -220
rect 732 -226 737 -206
rect 739 -213 744 -206
rect 782 -209 787 -206
rect 772 -212 777 -209
rect 739 -215 746 -213
rect 739 -217 742 -215
rect 744 -217 746 -215
rect 739 -219 746 -217
rect 750 -215 757 -212
rect 750 -217 752 -215
rect 754 -217 757 -215
rect 739 -226 744 -219
rect 750 -222 757 -217
rect 750 -224 752 -222
rect 754 -224 757 -222
rect 750 -226 757 -224
rect 759 -222 767 -212
rect 759 -224 762 -222
rect 764 -224 767 -222
rect 759 -226 767 -224
rect 769 -214 777 -212
rect 769 -216 772 -214
rect 774 -216 777 -214
rect 769 -219 777 -216
rect 779 -211 787 -209
rect 779 -213 782 -211
rect 784 -213 787 -211
rect 779 -219 787 -213
rect 789 -213 794 -206
rect 801 -209 807 -207
rect 801 -211 803 -209
rect 805 -211 807 -209
rect 801 -213 807 -211
rect 820 -209 826 -207
rect 867 -205 874 -203
rect 867 -207 870 -205
rect 872 -207 874 -205
rect 820 -211 822 -209
rect 824 -211 826 -209
rect 820 -213 826 -211
rect 789 -215 796 -213
rect 789 -217 792 -215
rect 794 -217 796 -215
rect 789 -219 796 -217
rect 769 -226 774 -219
rect 801 -220 806 -213
rect 822 -217 826 -213
rect 867 -213 874 -207
rect 849 -215 856 -213
rect 849 -217 851 -215
rect 853 -217 856 -215
rect 822 -220 828 -217
rect 801 -226 808 -220
rect 810 -222 818 -220
rect 810 -224 813 -222
rect 815 -224 818 -222
rect 810 -226 818 -224
rect 820 -226 828 -220
rect 830 -220 835 -217
rect 849 -219 856 -217
rect 830 -222 837 -220
rect 830 -224 833 -222
rect 835 -224 837 -222
rect 851 -224 856 -219
rect 858 -224 863 -213
rect 865 -215 874 -213
rect 891 -213 896 -206
rect 889 -215 896 -213
rect 865 -224 876 -215
rect 878 -217 885 -215
rect 878 -219 881 -217
rect 883 -219 885 -217
rect 889 -217 891 -215
rect 893 -217 896 -215
rect 889 -219 896 -217
rect 898 -209 903 -206
rect 898 -211 906 -209
rect 898 -213 901 -211
rect 903 -213 906 -211
rect 898 -219 906 -213
rect 908 -212 913 -209
rect 908 -214 916 -212
rect 908 -216 911 -214
rect 913 -216 916 -214
rect 908 -219 916 -216
rect 878 -221 885 -219
rect 878 -224 883 -221
rect 830 -226 837 -224
rect 911 -226 916 -219
rect 918 -222 926 -212
rect 918 -224 921 -222
rect 923 -224 926 -222
rect 918 -226 926 -224
rect 928 -215 935 -212
rect 941 -213 946 -206
rect 928 -217 931 -215
rect 933 -217 935 -215
rect 928 -222 935 -217
rect 939 -215 946 -213
rect 939 -217 941 -215
rect 943 -217 946 -215
rect 939 -219 946 -217
rect 928 -224 931 -222
rect 933 -224 935 -222
rect 928 -226 935 -224
rect 941 -226 946 -219
rect 948 -226 953 -206
rect 955 -208 964 -206
rect 955 -210 958 -208
rect 960 -210 964 -208
rect 955 -220 964 -210
rect 966 -213 971 -206
rect 981 -213 986 -206
rect 966 -215 973 -213
rect 966 -217 969 -215
rect 971 -217 973 -215
rect 966 -220 973 -217
rect 979 -215 986 -213
rect 979 -217 981 -215
rect 983 -217 986 -215
rect 979 -220 986 -217
rect 988 -208 997 -206
rect 988 -210 992 -208
rect 994 -210 997 -208
rect 988 -220 997 -210
rect 955 -226 962 -220
rect 990 -226 997 -220
rect 999 -226 1004 -206
rect 1006 -213 1011 -206
rect 1049 -209 1054 -206
rect 1039 -212 1044 -209
rect 1006 -215 1013 -213
rect 1006 -217 1009 -215
rect 1011 -217 1013 -215
rect 1006 -219 1013 -217
rect 1017 -215 1024 -212
rect 1017 -217 1019 -215
rect 1021 -217 1024 -215
rect 1006 -226 1011 -219
rect 1017 -222 1024 -217
rect 1017 -224 1019 -222
rect 1021 -224 1024 -222
rect 1017 -226 1024 -224
rect 1026 -222 1034 -212
rect 1026 -224 1029 -222
rect 1031 -224 1034 -222
rect 1026 -226 1034 -224
rect 1036 -214 1044 -212
rect 1036 -216 1039 -214
rect 1041 -216 1044 -214
rect 1036 -219 1044 -216
rect 1046 -211 1054 -209
rect 1046 -213 1049 -211
rect 1051 -213 1054 -211
rect 1046 -219 1054 -213
rect 1056 -213 1061 -206
rect 1068 -209 1074 -207
rect 1068 -211 1070 -209
rect 1072 -211 1074 -209
rect 1068 -213 1074 -211
rect 1087 -209 1093 -207
rect 1134 -205 1141 -203
rect 1134 -207 1137 -205
rect 1139 -207 1141 -205
rect 1087 -211 1089 -209
rect 1091 -211 1093 -209
rect 1087 -213 1093 -211
rect 1056 -215 1063 -213
rect 1056 -217 1059 -215
rect 1061 -217 1063 -215
rect 1056 -219 1063 -217
rect 1036 -226 1041 -219
rect 1068 -220 1073 -213
rect 1089 -217 1093 -213
rect 1134 -213 1141 -207
rect 1116 -215 1123 -213
rect 1116 -217 1118 -215
rect 1120 -217 1123 -215
rect 1089 -220 1095 -217
rect 1068 -226 1075 -220
rect 1077 -222 1085 -220
rect 1077 -224 1080 -222
rect 1082 -224 1085 -222
rect 1077 -226 1085 -224
rect 1087 -226 1095 -220
rect 1097 -220 1102 -217
rect 1116 -219 1123 -217
rect 1097 -222 1104 -220
rect 1097 -224 1100 -222
rect 1102 -224 1104 -222
rect 1118 -224 1123 -219
rect 1125 -224 1130 -213
rect 1132 -215 1141 -213
rect 1158 -213 1163 -206
rect 1156 -215 1163 -213
rect 1132 -224 1143 -215
rect 1145 -217 1152 -215
rect 1145 -219 1148 -217
rect 1150 -219 1152 -217
rect 1156 -217 1158 -215
rect 1160 -217 1163 -215
rect 1156 -219 1163 -217
rect 1165 -209 1170 -206
rect 1165 -211 1173 -209
rect 1165 -213 1168 -211
rect 1170 -213 1173 -211
rect 1165 -219 1173 -213
rect 1175 -212 1180 -209
rect 1175 -214 1183 -212
rect 1175 -216 1178 -214
rect 1180 -216 1183 -214
rect 1175 -219 1183 -216
rect 1145 -221 1152 -219
rect 1145 -224 1150 -221
rect 1097 -226 1104 -224
rect 1178 -226 1183 -219
rect 1185 -222 1193 -212
rect 1185 -224 1188 -222
rect 1190 -224 1193 -222
rect 1185 -226 1193 -224
rect 1195 -215 1202 -212
rect 1208 -213 1213 -206
rect 1195 -217 1198 -215
rect 1200 -217 1202 -215
rect 1195 -222 1202 -217
rect 1206 -215 1213 -213
rect 1206 -217 1208 -215
rect 1210 -217 1213 -215
rect 1206 -219 1213 -217
rect 1195 -224 1198 -222
rect 1200 -224 1202 -222
rect 1195 -226 1202 -224
rect 1208 -226 1213 -219
rect 1215 -226 1220 -206
rect 1222 -208 1231 -206
rect 1222 -210 1225 -208
rect 1227 -210 1231 -208
rect 1222 -220 1231 -210
rect 1233 -213 1238 -206
rect 1248 -213 1253 -206
rect 1233 -215 1240 -213
rect 1233 -217 1236 -215
rect 1238 -217 1240 -215
rect 1233 -220 1240 -217
rect 1246 -215 1253 -213
rect 1246 -217 1248 -215
rect 1250 -217 1253 -215
rect 1246 -220 1253 -217
rect 1255 -208 1264 -206
rect 1255 -210 1259 -208
rect 1261 -210 1264 -208
rect 1255 -220 1264 -210
rect 1222 -226 1229 -220
rect 1257 -226 1264 -220
rect 1266 -226 1271 -206
rect 1273 -213 1278 -206
rect 1316 -209 1321 -206
rect 1306 -212 1311 -209
rect 1273 -215 1280 -213
rect 1273 -217 1276 -215
rect 1278 -217 1280 -215
rect 1273 -219 1280 -217
rect 1284 -215 1291 -212
rect 1284 -217 1286 -215
rect 1288 -217 1291 -215
rect 1273 -226 1278 -219
rect 1284 -222 1291 -217
rect 1284 -224 1286 -222
rect 1288 -224 1291 -222
rect 1284 -226 1291 -224
rect 1293 -222 1301 -212
rect 1293 -224 1296 -222
rect 1298 -224 1301 -222
rect 1293 -226 1301 -224
rect 1303 -214 1311 -212
rect 1303 -216 1306 -214
rect 1308 -216 1311 -214
rect 1303 -219 1311 -216
rect 1313 -211 1321 -209
rect 1313 -213 1316 -211
rect 1318 -213 1321 -211
rect 1313 -219 1321 -213
rect 1323 -213 1328 -206
rect 1335 -209 1341 -207
rect 1335 -211 1337 -209
rect 1339 -211 1341 -209
rect 1335 -213 1341 -211
rect 1354 -209 1360 -207
rect 1401 -205 1408 -203
rect 1401 -207 1404 -205
rect 1406 -207 1408 -205
rect 1354 -211 1356 -209
rect 1358 -211 1360 -209
rect 1354 -213 1360 -211
rect 1323 -215 1330 -213
rect 1323 -217 1326 -215
rect 1328 -217 1330 -215
rect 1323 -219 1330 -217
rect 1303 -226 1308 -219
rect 1335 -220 1340 -213
rect 1356 -217 1360 -213
rect 1401 -213 1408 -207
rect 1383 -215 1390 -213
rect 1383 -217 1385 -215
rect 1387 -217 1390 -215
rect 1356 -220 1362 -217
rect 1335 -226 1342 -220
rect 1344 -222 1352 -220
rect 1344 -224 1347 -222
rect 1349 -224 1352 -222
rect 1344 -226 1352 -224
rect 1354 -226 1362 -220
rect 1364 -220 1369 -217
rect 1383 -219 1390 -217
rect 1364 -222 1371 -220
rect 1364 -224 1367 -222
rect 1369 -224 1371 -222
rect 1385 -224 1390 -219
rect 1392 -224 1397 -213
rect 1399 -215 1408 -213
rect 1425 -213 1430 -206
rect 1423 -215 1430 -213
rect 1399 -224 1410 -215
rect 1412 -217 1419 -215
rect 1412 -219 1415 -217
rect 1417 -219 1419 -217
rect 1423 -217 1425 -215
rect 1427 -217 1430 -215
rect 1423 -219 1430 -217
rect 1432 -209 1437 -206
rect 1432 -211 1440 -209
rect 1432 -213 1435 -211
rect 1437 -213 1440 -211
rect 1432 -219 1440 -213
rect 1442 -212 1447 -209
rect 1442 -214 1450 -212
rect 1442 -216 1445 -214
rect 1447 -216 1450 -214
rect 1442 -219 1450 -216
rect 1412 -221 1419 -219
rect 1412 -224 1417 -221
rect 1364 -226 1371 -224
rect 1445 -226 1450 -219
rect 1452 -222 1460 -212
rect 1452 -224 1455 -222
rect 1457 -224 1460 -222
rect 1452 -226 1460 -224
rect 1462 -215 1469 -212
rect 1475 -213 1480 -206
rect 1462 -217 1465 -215
rect 1467 -217 1469 -215
rect 1462 -222 1469 -217
rect 1473 -215 1480 -213
rect 1473 -217 1475 -215
rect 1477 -217 1480 -215
rect 1473 -219 1480 -217
rect 1462 -224 1465 -222
rect 1467 -224 1469 -222
rect 1462 -226 1469 -224
rect 1475 -226 1480 -219
rect 1482 -226 1487 -206
rect 1489 -208 1498 -206
rect 1489 -210 1492 -208
rect 1494 -210 1498 -208
rect 1489 -220 1498 -210
rect 1500 -213 1505 -206
rect 1515 -213 1520 -206
rect 1500 -215 1507 -213
rect 1500 -217 1503 -215
rect 1505 -217 1507 -215
rect 1500 -220 1507 -217
rect 1513 -215 1520 -213
rect 1513 -217 1515 -215
rect 1517 -217 1520 -215
rect 1513 -220 1520 -217
rect 1522 -208 1531 -206
rect 1522 -210 1526 -208
rect 1528 -210 1531 -208
rect 1522 -220 1531 -210
rect 1489 -226 1496 -220
rect 1524 -226 1531 -220
rect 1533 -226 1538 -206
rect 1540 -213 1545 -206
rect 1583 -209 1588 -206
rect 1573 -212 1578 -209
rect 1540 -215 1547 -213
rect 1540 -217 1543 -215
rect 1545 -217 1547 -215
rect 1540 -219 1547 -217
rect 1551 -215 1558 -212
rect 1551 -217 1553 -215
rect 1555 -217 1558 -215
rect 1540 -226 1545 -219
rect 1551 -222 1558 -217
rect 1551 -224 1553 -222
rect 1555 -224 1558 -222
rect 1551 -226 1558 -224
rect 1560 -222 1568 -212
rect 1560 -224 1563 -222
rect 1565 -224 1568 -222
rect 1560 -226 1568 -224
rect 1570 -214 1578 -212
rect 1570 -216 1573 -214
rect 1575 -216 1578 -214
rect 1570 -219 1578 -216
rect 1580 -211 1588 -209
rect 1580 -213 1583 -211
rect 1585 -213 1588 -211
rect 1580 -219 1588 -213
rect 1590 -213 1595 -206
rect 1602 -209 1608 -207
rect 1602 -211 1604 -209
rect 1606 -211 1608 -209
rect 1602 -213 1608 -211
rect 1621 -209 1627 -207
rect 1668 -205 1675 -203
rect 1668 -207 1671 -205
rect 1673 -207 1675 -205
rect 1621 -211 1623 -209
rect 1625 -211 1627 -209
rect 1621 -213 1627 -211
rect 1590 -215 1597 -213
rect 1590 -217 1593 -215
rect 1595 -217 1597 -215
rect 1590 -219 1597 -217
rect 1570 -226 1575 -219
rect 1602 -220 1607 -213
rect 1623 -217 1627 -213
rect 1668 -213 1675 -207
rect 1650 -215 1657 -213
rect 1650 -217 1652 -215
rect 1654 -217 1657 -215
rect 1623 -220 1629 -217
rect 1602 -226 1609 -220
rect 1611 -222 1619 -220
rect 1611 -224 1614 -222
rect 1616 -224 1619 -222
rect 1611 -226 1619 -224
rect 1621 -226 1629 -220
rect 1631 -220 1636 -217
rect 1650 -219 1657 -217
rect 1631 -222 1638 -220
rect 1631 -224 1634 -222
rect 1636 -224 1638 -222
rect 1652 -224 1657 -219
rect 1659 -224 1664 -213
rect 1666 -215 1675 -213
rect 1692 -213 1697 -206
rect 1690 -215 1697 -213
rect 1666 -224 1677 -215
rect 1679 -217 1686 -215
rect 1679 -219 1682 -217
rect 1684 -219 1686 -217
rect 1690 -217 1692 -215
rect 1694 -217 1697 -215
rect 1690 -219 1697 -217
rect 1699 -209 1704 -206
rect 1699 -211 1707 -209
rect 1699 -213 1702 -211
rect 1704 -213 1707 -211
rect 1699 -219 1707 -213
rect 1709 -212 1714 -209
rect 1709 -214 1717 -212
rect 1709 -216 1712 -214
rect 1714 -216 1717 -214
rect 1709 -219 1717 -216
rect 1679 -221 1686 -219
rect 1679 -224 1684 -221
rect 1631 -226 1638 -224
rect 1712 -226 1717 -219
rect 1719 -222 1727 -212
rect 1719 -224 1722 -222
rect 1724 -224 1727 -222
rect 1719 -226 1727 -224
rect 1729 -215 1736 -212
rect 1742 -213 1747 -206
rect 1729 -217 1732 -215
rect 1734 -217 1736 -215
rect 1729 -222 1736 -217
rect 1740 -215 1747 -213
rect 1740 -217 1742 -215
rect 1744 -217 1747 -215
rect 1740 -219 1747 -217
rect 1729 -224 1732 -222
rect 1734 -224 1736 -222
rect 1729 -226 1736 -224
rect 1742 -226 1747 -219
rect 1749 -226 1754 -206
rect 1756 -208 1765 -206
rect 1756 -210 1759 -208
rect 1761 -210 1765 -208
rect 1756 -220 1765 -210
rect 1767 -213 1772 -206
rect 1782 -213 1787 -206
rect 1767 -215 1774 -213
rect 1767 -217 1770 -215
rect 1772 -217 1774 -215
rect 1767 -220 1774 -217
rect 1780 -215 1787 -213
rect 1780 -217 1782 -215
rect 1784 -217 1787 -215
rect 1780 -220 1787 -217
rect 1789 -208 1798 -206
rect 1789 -210 1793 -208
rect 1795 -210 1798 -208
rect 1789 -220 1798 -210
rect 1756 -226 1763 -220
rect 1791 -226 1798 -220
rect 1800 -226 1805 -206
rect 1807 -213 1812 -206
rect 1850 -209 1855 -206
rect 1840 -212 1845 -209
rect 1807 -215 1814 -213
rect 1807 -217 1810 -215
rect 1812 -217 1814 -215
rect 1807 -219 1814 -217
rect 1818 -215 1825 -212
rect 1818 -217 1820 -215
rect 1822 -217 1825 -215
rect 1807 -226 1812 -219
rect 1818 -222 1825 -217
rect 1818 -224 1820 -222
rect 1822 -224 1825 -222
rect 1818 -226 1825 -224
rect 1827 -222 1835 -212
rect 1827 -224 1830 -222
rect 1832 -224 1835 -222
rect 1827 -226 1835 -224
rect 1837 -214 1845 -212
rect 1837 -216 1840 -214
rect 1842 -216 1845 -214
rect 1837 -219 1845 -216
rect 1847 -211 1855 -209
rect 1847 -213 1850 -211
rect 1852 -213 1855 -211
rect 1847 -219 1855 -213
rect 1857 -213 1862 -206
rect 1869 -209 1875 -207
rect 1869 -211 1871 -209
rect 1873 -211 1875 -209
rect 1869 -213 1875 -211
rect 1888 -209 1894 -207
rect 1888 -211 1890 -209
rect 1892 -211 1894 -209
rect 1888 -213 1894 -211
rect 1966 -205 1972 -203
rect 1966 -207 1968 -205
rect 1970 -207 1972 -205
rect 1966 -209 1972 -207
rect 1950 -212 1955 -209
rect 1857 -215 1864 -213
rect 1857 -217 1860 -215
rect 1862 -217 1864 -215
rect 1857 -219 1864 -217
rect 1837 -226 1842 -219
rect 1869 -220 1874 -213
rect 1890 -217 1894 -213
rect 1926 -214 1935 -212
rect 1926 -216 1928 -214
rect 1930 -216 1935 -214
rect 1926 -217 1935 -216
rect 1890 -220 1896 -217
rect 1869 -226 1876 -220
rect 1878 -222 1886 -220
rect 1878 -224 1881 -222
rect 1883 -224 1886 -222
rect 1878 -226 1886 -224
rect 1888 -226 1896 -220
rect 1898 -220 1903 -217
rect 1914 -220 1919 -217
rect 1898 -222 1905 -220
rect 1898 -224 1901 -222
rect 1903 -224 1905 -222
rect 1898 -226 1905 -224
rect 1912 -222 1919 -220
rect 1912 -224 1914 -222
rect 1916 -224 1919 -222
rect 1912 -226 1919 -224
rect 1921 -221 1935 -217
rect 1937 -217 1945 -212
rect 1937 -219 1940 -217
rect 1942 -219 1945 -217
rect 1937 -221 1945 -219
rect 1947 -215 1955 -212
rect 1947 -217 1950 -215
rect 1952 -217 1955 -215
rect 1947 -221 1955 -217
rect 1957 -221 1962 -209
rect 1964 -221 1972 -209
rect 1978 -213 1983 -206
rect 1976 -215 1983 -213
rect 1976 -217 1978 -215
rect 1980 -217 1983 -215
rect 1976 -219 1983 -217
rect 1985 -209 1990 -206
rect 1985 -211 1993 -209
rect 1985 -213 1988 -211
rect 1990 -213 1993 -211
rect 1985 -219 1993 -213
rect 1995 -212 2000 -209
rect 1995 -214 2003 -212
rect 1995 -216 1998 -214
rect 2000 -216 2003 -214
rect 1995 -219 2003 -216
rect 1921 -226 1926 -221
rect 1998 -226 2003 -219
rect 2005 -222 2013 -212
rect 2005 -224 2008 -222
rect 2010 -224 2013 -222
rect 2005 -226 2013 -224
rect 2015 -215 2022 -212
rect 2028 -213 2033 -206
rect 2015 -217 2018 -215
rect 2020 -217 2022 -215
rect 2015 -222 2022 -217
rect 2026 -215 2033 -213
rect 2026 -217 2028 -215
rect 2030 -217 2033 -215
rect 2026 -219 2033 -217
rect 2015 -224 2018 -222
rect 2020 -224 2022 -222
rect 2015 -226 2022 -224
rect 2028 -226 2033 -219
rect 2035 -226 2040 -206
rect 2042 -208 2051 -206
rect 2042 -210 2045 -208
rect 2047 -210 2051 -208
rect 2042 -220 2051 -210
rect 2053 -213 2058 -206
rect 2068 -213 2073 -206
rect 2053 -215 2060 -213
rect 2053 -217 2056 -215
rect 2058 -217 2060 -215
rect 2053 -220 2060 -217
rect 2066 -215 2073 -213
rect 2066 -217 2068 -215
rect 2070 -217 2073 -215
rect 2066 -220 2073 -217
rect 2075 -208 2084 -206
rect 2075 -210 2079 -208
rect 2081 -210 2084 -208
rect 2075 -220 2084 -210
rect 2042 -226 2049 -220
rect 2077 -226 2084 -220
rect 2086 -226 2091 -206
rect 2093 -213 2098 -206
rect 2136 -209 2141 -206
rect 2126 -212 2131 -209
rect 2093 -215 2100 -213
rect 2093 -217 2096 -215
rect 2098 -217 2100 -215
rect 2093 -219 2100 -217
rect 2104 -215 2111 -212
rect 2104 -217 2106 -215
rect 2108 -217 2111 -215
rect 2093 -226 2098 -219
rect 2104 -222 2111 -217
rect 2104 -224 2106 -222
rect 2108 -224 2111 -222
rect 2104 -226 2111 -224
rect 2113 -222 2121 -212
rect 2113 -224 2116 -222
rect 2118 -224 2121 -222
rect 2113 -226 2121 -224
rect 2123 -214 2131 -212
rect 2123 -216 2126 -214
rect 2128 -216 2131 -214
rect 2123 -219 2131 -216
rect 2133 -211 2141 -209
rect 2133 -213 2136 -211
rect 2138 -213 2141 -211
rect 2133 -219 2141 -213
rect 2143 -213 2148 -206
rect 2155 -209 2161 -207
rect 2155 -211 2157 -209
rect 2159 -211 2161 -209
rect 2155 -213 2161 -211
rect 2174 -209 2180 -207
rect 2174 -211 2176 -209
rect 2178 -211 2180 -209
rect 2174 -213 2180 -211
rect 2143 -215 2150 -213
rect 2143 -217 2146 -215
rect 2148 -217 2150 -215
rect 2143 -219 2150 -217
rect 2123 -226 2128 -219
rect 2155 -220 2160 -213
rect 2176 -217 2180 -213
rect 2210 -214 2216 -212
rect 2199 -216 2206 -214
rect 2176 -220 2182 -217
rect 2155 -226 2162 -220
rect 2164 -222 2172 -220
rect 2164 -224 2167 -222
rect 2169 -224 2172 -222
rect 2164 -226 2172 -224
rect 2174 -226 2182 -220
rect 2184 -220 2189 -217
rect 2199 -218 2201 -216
rect 2203 -218 2206 -216
rect 2199 -220 2206 -218
rect 2208 -216 2216 -214
rect 2208 -218 2211 -216
rect 2213 -218 2216 -216
rect 2208 -220 2216 -218
rect 2218 -220 2223 -212
rect 2225 -214 2233 -212
rect 2225 -216 2228 -214
rect 2230 -216 2233 -214
rect 2225 -220 2233 -216
rect 2235 -220 2240 -212
rect 2242 -214 2250 -212
rect 2242 -216 2245 -214
rect 2247 -216 2250 -214
rect 2242 -220 2250 -216
rect 2184 -222 2191 -220
rect 2184 -224 2187 -222
rect 2189 -224 2191 -222
rect 2184 -226 2191 -224
rect 2245 -221 2250 -220
rect 2252 -215 2257 -212
rect 2278 -214 2284 -212
rect 2252 -217 2259 -215
rect 2252 -219 2255 -217
rect 2257 -219 2259 -217
rect 2252 -221 2259 -219
rect 2267 -216 2274 -214
rect 2267 -218 2269 -216
rect 2271 -218 2274 -216
rect 2267 -220 2274 -218
rect 2276 -216 2284 -214
rect 2276 -218 2279 -216
rect 2281 -218 2284 -216
rect 2276 -220 2284 -218
rect 2286 -220 2291 -212
rect 2293 -214 2301 -212
rect 2293 -216 2296 -214
rect 2298 -216 2301 -214
rect 2293 -220 2301 -216
rect 2303 -220 2308 -212
rect 2310 -214 2318 -212
rect 2310 -216 2313 -214
rect 2315 -216 2318 -214
rect 2310 -220 2318 -216
rect 2313 -221 2318 -220
rect 2320 -215 2325 -212
rect 2320 -217 2327 -215
rect 2320 -219 2323 -217
rect 2325 -219 2327 -217
rect 2320 -221 2327 -219
<< pdif >>
rect 8 289 15 291
rect 8 287 10 289
rect 12 287 15 289
rect 8 278 15 287
rect 17 289 25 291
rect 17 287 20 289
rect 22 287 25 289
rect 17 282 25 287
rect 17 280 20 282
rect 22 280 25 282
rect 17 278 25 280
rect 27 289 33 291
rect 48 289 55 291
rect 27 287 35 289
rect 27 285 30 287
rect 32 285 35 287
rect 27 278 35 285
rect 29 271 35 278
rect 37 284 42 289
rect 48 287 50 289
rect 52 287 55 289
rect 37 282 44 284
rect 37 280 40 282
rect 42 280 44 282
rect 37 275 44 280
rect 48 278 55 287
rect 57 289 65 291
rect 57 287 60 289
rect 62 287 65 289
rect 57 282 65 287
rect 57 280 60 282
rect 62 280 65 282
rect 57 278 65 280
rect 67 289 73 291
rect 67 287 75 289
rect 67 285 70 287
rect 72 285 75 287
rect 67 278 75 285
rect 37 273 40 275
rect 42 273 44 275
rect 37 271 44 273
rect 69 271 75 278
rect 77 284 82 289
rect 90 286 95 298
rect 88 284 95 286
rect 77 282 84 284
rect 77 280 80 282
rect 82 280 84 282
rect 77 275 84 280
rect 77 273 80 275
rect 82 273 84 275
rect 88 282 90 284
rect 92 282 95 284
rect 88 277 95 282
rect 88 275 90 277
rect 92 275 95 277
rect 88 273 95 275
rect 97 296 106 298
rect 97 294 101 296
rect 103 294 106 296
rect 129 296 143 298
rect 129 295 136 296
rect 97 286 106 294
rect 113 286 118 295
rect 97 273 108 286
rect 110 277 118 286
rect 110 275 113 277
rect 115 275 118 277
rect 110 273 118 275
rect 77 271 84 273
rect 113 270 118 273
rect 120 270 125 295
rect 127 294 136 295
rect 138 294 143 296
rect 127 289 143 294
rect 127 287 136 289
rect 138 287 143 289
rect 127 270 143 287
rect 145 288 153 298
rect 145 286 148 288
rect 150 286 153 288
rect 145 281 153 286
rect 145 279 148 281
rect 150 279 153 281
rect 145 270 153 279
rect 155 296 163 298
rect 155 294 158 296
rect 160 294 163 296
rect 155 289 163 294
rect 155 287 158 289
rect 160 287 163 289
rect 155 270 163 287
rect 165 283 170 298
rect 180 283 185 298
rect 165 281 172 283
rect 165 279 168 281
rect 170 279 172 281
rect 165 274 172 279
rect 165 272 168 274
rect 170 272 172 274
rect 165 270 172 272
rect 178 281 185 283
rect 178 279 180 281
rect 182 279 185 281
rect 178 274 185 279
rect 178 272 180 274
rect 182 272 185 274
rect 178 270 185 272
rect 187 296 195 298
rect 187 294 190 296
rect 192 294 195 296
rect 187 289 195 294
rect 187 287 190 289
rect 192 287 195 289
rect 187 270 195 287
rect 197 288 205 298
rect 197 286 200 288
rect 202 286 205 288
rect 197 281 205 286
rect 197 279 200 281
rect 202 279 205 281
rect 197 270 205 279
rect 207 296 221 298
rect 207 294 212 296
rect 214 295 221 296
rect 244 296 253 298
rect 214 294 223 295
rect 207 289 223 294
rect 207 287 212 289
rect 214 287 223 289
rect 207 270 223 287
rect 225 270 230 295
rect 232 286 237 295
rect 244 294 247 296
rect 249 294 253 296
rect 244 286 253 294
rect 232 277 240 286
rect 232 275 235 277
rect 237 275 240 277
rect 232 273 240 275
rect 242 273 253 286
rect 255 286 260 298
rect 269 291 274 298
rect 267 289 274 291
rect 267 287 269 289
rect 271 287 274 289
rect 255 284 262 286
rect 267 285 274 287
rect 255 282 258 284
rect 260 282 262 284
rect 255 277 262 282
rect 269 277 274 285
rect 276 277 281 298
rect 283 296 292 298
rect 283 294 288 296
rect 290 294 292 296
rect 283 288 292 294
rect 315 289 322 291
rect 283 277 294 288
rect 255 275 258 277
rect 260 275 262 277
rect 255 273 262 275
rect 232 270 237 273
rect 286 270 294 277
rect 296 286 303 288
rect 296 284 299 286
rect 301 284 303 286
rect 296 279 303 284
rect 296 277 299 279
rect 301 277 303 279
rect 315 287 317 289
rect 319 287 322 289
rect 315 278 322 287
rect 324 289 332 291
rect 324 287 327 289
rect 329 287 332 289
rect 324 282 332 287
rect 324 280 327 282
rect 329 280 332 282
rect 324 278 332 280
rect 334 289 340 291
rect 334 287 342 289
rect 334 285 337 287
rect 339 285 342 287
rect 334 278 342 285
rect 296 275 303 277
rect 296 270 301 275
rect 336 271 342 278
rect 344 284 349 289
rect 357 286 362 298
rect 355 284 362 286
rect 344 282 351 284
rect 344 280 347 282
rect 349 280 351 282
rect 344 275 351 280
rect 344 273 347 275
rect 349 273 351 275
rect 355 282 357 284
rect 359 282 362 284
rect 355 277 362 282
rect 355 275 357 277
rect 359 275 362 277
rect 355 273 362 275
rect 364 296 373 298
rect 364 294 368 296
rect 370 294 373 296
rect 396 296 410 298
rect 396 295 403 296
rect 364 286 373 294
rect 380 286 385 295
rect 364 273 375 286
rect 377 277 385 286
rect 377 275 380 277
rect 382 275 385 277
rect 377 273 385 275
rect 344 271 351 273
rect 380 270 385 273
rect 387 270 392 295
rect 394 294 403 295
rect 405 294 410 296
rect 394 289 410 294
rect 394 287 403 289
rect 405 287 410 289
rect 394 270 410 287
rect 412 288 420 298
rect 412 286 415 288
rect 417 286 420 288
rect 412 281 420 286
rect 412 279 415 281
rect 417 279 420 281
rect 412 270 420 279
rect 422 296 430 298
rect 422 294 425 296
rect 427 294 430 296
rect 422 289 430 294
rect 422 287 425 289
rect 427 287 430 289
rect 422 270 430 287
rect 432 283 437 298
rect 447 283 452 298
rect 432 281 439 283
rect 432 279 435 281
rect 437 279 439 281
rect 432 274 439 279
rect 432 272 435 274
rect 437 272 439 274
rect 432 270 439 272
rect 445 281 452 283
rect 445 279 447 281
rect 449 279 452 281
rect 445 274 452 279
rect 445 272 447 274
rect 449 272 452 274
rect 445 270 452 272
rect 454 296 462 298
rect 454 294 457 296
rect 459 294 462 296
rect 454 289 462 294
rect 454 287 457 289
rect 459 287 462 289
rect 454 270 462 287
rect 464 288 472 298
rect 464 286 467 288
rect 469 286 472 288
rect 464 281 472 286
rect 464 279 467 281
rect 469 279 472 281
rect 464 270 472 279
rect 474 296 488 298
rect 474 294 479 296
rect 481 295 488 296
rect 511 296 520 298
rect 481 294 490 295
rect 474 289 490 294
rect 474 287 479 289
rect 481 287 490 289
rect 474 270 490 287
rect 492 270 497 295
rect 499 286 504 295
rect 511 294 514 296
rect 516 294 520 296
rect 511 286 520 294
rect 499 277 507 286
rect 499 275 502 277
rect 504 275 507 277
rect 499 273 507 275
rect 509 273 520 286
rect 522 286 527 298
rect 536 291 541 298
rect 534 289 541 291
rect 534 287 536 289
rect 538 287 541 289
rect 522 284 529 286
rect 534 285 541 287
rect 522 282 525 284
rect 527 282 529 284
rect 522 277 529 282
rect 536 277 541 285
rect 543 277 548 298
rect 550 296 559 298
rect 550 294 555 296
rect 557 294 559 296
rect 550 288 559 294
rect 582 289 589 291
rect 550 277 561 288
rect 522 275 525 277
rect 527 275 529 277
rect 522 273 529 275
rect 499 270 504 273
rect 553 270 561 277
rect 563 286 570 288
rect 563 284 566 286
rect 568 284 570 286
rect 563 279 570 284
rect 563 277 566 279
rect 568 277 570 279
rect 582 287 584 289
rect 586 287 589 289
rect 582 278 589 287
rect 591 289 599 291
rect 591 287 594 289
rect 596 287 599 289
rect 591 282 599 287
rect 591 280 594 282
rect 596 280 599 282
rect 591 278 599 280
rect 601 289 607 291
rect 601 287 609 289
rect 601 285 604 287
rect 606 285 609 287
rect 601 278 609 285
rect 563 275 570 277
rect 563 270 568 275
rect 603 271 609 278
rect 611 284 616 289
rect 624 286 629 298
rect 622 284 629 286
rect 611 282 618 284
rect 611 280 614 282
rect 616 280 618 282
rect 611 275 618 280
rect 611 273 614 275
rect 616 273 618 275
rect 622 282 624 284
rect 626 282 629 284
rect 622 277 629 282
rect 622 275 624 277
rect 626 275 629 277
rect 622 273 629 275
rect 631 296 640 298
rect 631 294 635 296
rect 637 294 640 296
rect 663 296 677 298
rect 663 295 670 296
rect 631 286 640 294
rect 647 286 652 295
rect 631 273 642 286
rect 644 277 652 286
rect 644 275 647 277
rect 649 275 652 277
rect 644 273 652 275
rect 611 271 618 273
rect 647 270 652 273
rect 654 270 659 295
rect 661 294 670 295
rect 672 294 677 296
rect 661 289 677 294
rect 661 287 670 289
rect 672 287 677 289
rect 661 270 677 287
rect 679 288 687 298
rect 679 286 682 288
rect 684 286 687 288
rect 679 281 687 286
rect 679 279 682 281
rect 684 279 687 281
rect 679 270 687 279
rect 689 296 697 298
rect 689 294 692 296
rect 694 294 697 296
rect 689 289 697 294
rect 689 287 692 289
rect 694 287 697 289
rect 689 270 697 287
rect 699 283 704 298
rect 714 283 719 298
rect 699 281 706 283
rect 699 279 702 281
rect 704 279 706 281
rect 699 274 706 279
rect 699 272 702 274
rect 704 272 706 274
rect 699 270 706 272
rect 712 281 719 283
rect 712 279 714 281
rect 716 279 719 281
rect 712 274 719 279
rect 712 272 714 274
rect 716 272 719 274
rect 712 270 719 272
rect 721 296 729 298
rect 721 294 724 296
rect 726 294 729 296
rect 721 289 729 294
rect 721 287 724 289
rect 726 287 729 289
rect 721 270 729 287
rect 731 288 739 298
rect 731 286 734 288
rect 736 286 739 288
rect 731 281 739 286
rect 731 279 734 281
rect 736 279 739 281
rect 731 270 739 279
rect 741 296 755 298
rect 741 294 746 296
rect 748 295 755 296
rect 778 296 787 298
rect 748 294 757 295
rect 741 289 757 294
rect 741 287 746 289
rect 748 287 757 289
rect 741 270 757 287
rect 759 270 764 295
rect 766 286 771 295
rect 778 294 781 296
rect 783 294 787 296
rect 778 286 787 294
rect 766 277 774 286
rect 766 275 769 277
rect 771 275 774 277
rect 766 273 774 275
rect 776 273 787 286
rect 789 286 794 298
rect 803 291 808 298
rect 801 289 808 291
rect 801 287 803 289
rect 805 287 808 289
rect 789 284 796 286
rect 801 285 808 287
rect 789 282 792 284
rect 794 282 796 284
rect 789 277 796 282
rect 803 277 808 285
rect 810 277 815 298
rect 817 296 826 298
rect 817 294 822 296
rect 824 294 826 296
rect 817 288 826 294
rect 849 289 856 291
rect 817 277 828 288
rect 789 275 792 277
rect 794 275 796 277
rect 789 273 796 275
rect 766 270 771 273
rect 820 270 828 277
rect 830 286 837 288
rect 830 284 833 286
rect 835 284 837 286
rect 830 279 837 284
rect 830 277 833 279
rect 835 277 837 279
rect 849 287 851 289
rect 853 287 856 289
rect 849 278 856 287
rect 858 289 866 291
rect 858 287 861 289
rect 863 287 866 289
rect 858 282 866 287
rect 858 280 861 282
rect 863 280 866 282
rect 858 278 866 280
rect 868 289 874 291
rect 868 287 876 289
rect 868 285 871 287
rect 873 285 876 287
rect 868 278 876 285
rect 830 275 837 277
rect 830 270 835 275
rect 870 271 876 278
rect 878 284 883 289
rect 891 286 896 298
rect 889 284 896 286
rect 878 282 885 284
rect 878 280 881 282
rect 883 280 885 282
rect 878 275 885 280
rect 878 273 881 275
rect 883 273 885 275
rect 889 282 891 284
rect 893 282 896 284
rect 889 277 896 282
rect 889 275 891 277
rect 893 275 896 277
rect 889 273 896 275
rect 898 296 907 298
rect 898 294 902 296
rect 904 294 907 296
rect 930 296 944 298
rect 930 295 937 296
rect 898 286 907 294
rect 914 286 919 295
rect 898 273 909 286
rect 911 277 919 286
rect 911 275 914 277
rect 916 275 919 277
rect 911 273 919 275
rect 878 271 885 273
rect 914 270 919 273
rect 921 270 926 295
rect 928 294 937 295
rect 939 294 944 296
rect 928 289 944 294
rect 928 287 937 289
rect 939 287 944 289
rect 928 270 944 287
rect 946 288 954 298
rect 946 286 949 288
rect 951 286 954 288
rect 946 281 954 286
rect 946 279 949 281
rect 951 279 954 281
rect 946 270 954 279
rect 956 296 964 298
rect 956 294 959 296
rect 961 294 964 296
rect 956 289 964 294
rect 956 287 959 289
rect 961 287 964 289
rect 956 270 964 287
rect 966 283 971 298
rect 981 283 986 298
rect 966 281 973 283
rect 966 279 969 281
rect 971 279 973 281
rect 966 274 973 279
rect 966 272 969 274
rect 971 272 973 274
rect 966 270 973 272
rect 979 281 986 283
rect 979 279 981 281
rect 983 279 986 281
rect 979 274 986 279
rect 979 272 981 274
rect 983 272 986 274
rect 979 270 986 272
rect 988 296 996 298
rect 988 294 991 296
rect 993 294 996 296
rect 988 289 996 294
rect 988 287 991 289
rect 993 287 996 289
rect 988 270 996 287
rect 998 288 1006 298
rect 998 286 1001 288
rect 1003 286 1006 288
rect 998 281 1006 286
rect 998 279 1001 281
rect 1003 279 1006 281
rect 998 270 1006 279
rect 1008 296 1022 298
rect 1008 294 1013 296
rect 1015 295 1022 296
rect 1045 296 1054 298
rect 1015 294 1024 295
rect 1008 289 1024 294
rect 1008 287 1013 289
rect 1015 287 1024 289
rect 1008 270 1024 287
rect 1026 270 1031 295
rect 1033 286 1038 295
rect 1045 294 1048 296
rect 1050 294 1054 296
rect 1045 286 1054 294
rect 1033 277 1041 286
rect 1033 275 1036 277
rect 1038 275 1041 277
rect 1033 273 1041 275
rect 1043 273 1054 286
rect 1056 286 1061 298
rect 1070 291 1075 298
rect 1068 289 1075 291
rect 1068 287 1070 289
rect 1072 287 1075 289
rect 1056 284 1063 286
rect 1068 285 1075 287
rect 1056 282 1059 284
rect 1061 282 1063 284
rect 1056 277 1063 282
rect 1070 277 1075 285
rect 1077 277 1082 298
rect 1084 296 1093 298
rect 1084 294 1089 296
rect 1091 294 1093 296
rect 1084 288 1093 294
rect 1116 289 1123 291
rect 1084 277 1095 288
rect 1056 275 1059 277
rect 1061 275 1063 277
rect 1056 273 1063 275
rect 1033 270 1038 273
rect 1087 270 1095 277
rect 1097 286 1104 288
rect 1097 284 1100 286
rect 1102 284 1104 286
rect 1097 279 1104 284
rect 1097 277 1100 279
rect 1102 277 1104 279
rect 1116 287 1118 289
rect 1120 287 1123 289
rect 1116 278 1123 287
rect 1125 289 1133 291
rect 1125 287 1128 289
rect 1130 287 1133 289
rect 1125 282 1133 287
rect 1125 280 1128 282
rect 1130 280 1133 282
rect 1125 278 1133 280
rect 1135 289 1141 291
rect 1135 287 1143 289
rect 1135 285 1138 287
rect 1140 285 1143 287
rect 1135 278 1143 285
rect 1097 275 1104 277
rect 1097 270 1102 275
rect 1137 271 1143 278
rect 1145 284 1150 289
rect 1158 286 1163 298
rect 1156 284 1163 286
rect 1145 282 1152 284
rect 1145 280 1148 282
rect 1150 280 1152 282
rect 1145 275 1152 280
rect 1145 273 1148 275
rect 1150 273 1152 275
rect 1156 282 1158 284
rect 1160 282 1163 284
rect 1156 277 1163 282
rect 1156 275 1158 277
rect 1160 275 1163 277
rect 1156 273 1163 275
rect 1165 296 1174 298
rect 1165 294 1169 296
rect 1171 294 1174 296
rect 1197 296 1211 298
rect 1197 295 1204 296
rect 1165 286 1174 294
rect 1181 286 1186 295
rect 1165 273 1176 286
rect 1178 277 1186 286
rect 1178 275 1181 277
rect 1183 275 1186 277
rect 1178 273 1186 275
rect 1145 271 1152 273
rect 1181 270 1186 273
rect 1188 270 1193 295
rect 1195 294 1204 295
rect 1206 294 1211 296
rect 1195 289 1211 294
rect 1195 287 1204 289
rect 1206 287 1211 289
rect 1195 270 1211 287
rect 1213 288 1221 298
rect 1213 286 1216 288
rect 1218 286 1221 288
rect 1213 281 1221 286
rect 1213 279 1216 281
rect 1218 279 1221 281
rect 1213 270 1221 279
rect 1223 296 1231 298
rect 1223 294 1226 296
rect 1228 294 1231 296
rect 1223 289 1231 294
rect 1223 287 1226 289
rect 1228 287 1231 289
rect 1223 270 1231 287
rect 1233 283 1238 298
rect 1248 283 1253 298
rect 1233 281 1240 283
rect 1233 279 1236 281
rect 1238 279 1240 281
rect 1233 274 1240 279
rect 1233 272 1236 274
rect 1238 272 1240 274
rect 1233 270 1240 272
rect 1246 281 1253 283
rect 1246 279 1248 281
rect 1250 279 1253 281
rect 1246 274 1253 279
rect 1246 272 1248 274
rect 1250 272 1253 274
rect 1246 270 1253 272
rect 1255 296 1263 298
rect 1255 294 1258 296
rect 1260 294 1263 296
rect 1255 289 1263 294
rect 1255 287 1258 289
rect 1260 287 1263 289
rect 1255 270 1263 287
rect 1265 288 1273 298
rect 1265 286 1268 288
rect 1270 286 1273 288
rect 1265 281 1273 286
rect 1265 279 1268 281
rect 1270 279 1273 281
rect 1265 270 1273 279
rect 1275 296 1289 298
rect 1275 294 1280 296
rect 1282 295 1289 296
rect 1312 296 1321 298
rect 1282 294 1291 295
rect 1275 289 1291 294
rect 1275 287 1280 289
rect 1282 287 1291 289
rect 1275 270 1291 287
rect 1293 270 1298 295
rect 1300 286 1305 295
rect 1312 294 1315 296
rect 1317 294 1321 296
rect 1312 286 1321 294
rect 1300 277 1308 286
rect 1300 275 1303 277
rect 1305 275 1308 277
rect 1300 273 1308 275
rect 1310 273 1321 286
rect 1323 286 1328 298
rect 1337 291 1342 298
rect 1335 289 1342 291
rect 1335 287 1337 289
rect 1339 287 1342 289
rect 1323 284 1330 286
rect 1335 285 1342 287
rect 1323 282 1326 284
rect 1328 282 1330 284
rect 1323 277 1330 282
rect 1337 277 1342 285
rect 1344 277 1349 298
rect 1351 296 1360 298
rect 1351 294 1356 296
rect 1358 294 1360 296
rect 1351 288 1360 294
rect 1383 289 1390 291
rect 1351 277 1362 288
rect 1323 275 1326 277
rect 1328 275 1330 277
rect 1323 273 1330 275
rect 1300 270 1305 273
rect 1354 270 1362 277
rect 1364 286 1371 288
rect 1364 284 1367 286
rect 1369 284 1371 286
rect 1364 279 1371 284
rect 1364 277 1367 279
rect 1369 277 1371 279
rect 1383 287 1385 289
rect 1387 287 1390 289
rect 1383 278 1390 287
rect 1392 289 1400 291
rect 1392 287 1395 289
rect 1397 287 1400 289
rect 1392 282 1400 287
rect 1392 280 1395 282
rect 1397 280 1400 282
rect 1392 278 1400 280
rect 1402 289 1408 291
rect 1402 287 1410 289
rect 1402 285 1405 287
rect 1407 285 1410 287
rect 1402 278 1410 285
rect 1364 275 1371 277
rect 1364 270 1369 275
rect 1404 271 1410 278
rect 1412 284 1417 289
rect 1425 286 1430 298
rect 1423 284 1430 286
rect 1412 282 1419 284
rect 1412 280 1415 282
rect 1417 280 1419 282
rect 1412 275 1419 280
rect 1412 273 1415 275
rect 1417 273 1419 275
rect 1423 282 1425 284
rect 1427 282 1430 284
rect 1423 277 1430 282
rect 1423 275 1425 277
rect 1427 275 1430 277
rect 1423 273 1430 275
rect 1432 296 1441 298
rect 1432 294 1436 296
rect 1438 294 1441 296
rect 1464 296 1478 298
rect 1464 295 1471 296
rect 1432 286 1441 294
rect 1448 286 1453 295
rect 1432 273 1443 286
rect 1445 277 1453 286
rect 1445 275 1448 277
rect 1450 275 1453 277
rect 1445 273 1453 275
rect 1412 271 1419 273
rect 1448 270 1453 273
rect 1455 270 1460 295
rect 1462 294 1471 295
rect 1473 294 1478 296
rect 1462 289 1478 294
rect 1462 287 1471 289
rect 1473 287 1478 289
rect 1462 270 1478 287
rect 1480 288 1488 298
rect 1480 286 1483 288
rect 1485 286 1488 288
rect 1480 281 1488 286
rect 1480 279 1483 281
rect 1485 279 1488 281
rect 1480 270 1488 279
rect 1490 296 1498 298
rect 1490 294 1493 296
rect 1495 294 1498 296
rect 1490 289 1498 294
rect 1490 287 1493 289
rect 1495 287 1498 289
rect 1490 270 1498 287
rect 1500 283 1505 298
rect 1515 283 1520 298
rect 1500 281 1507 283
rect 1500 279 1503 281
rect 1505 279 1507 281
rect 1500 274 1507 279
rect 1500 272 1503 274
rect 1505 272 1507 274
rect 1500 270 1507 272
rect 1513 281 1520 283
rect 1513 279 1515 281
rect 1517 279 1520 281
rect 1513 274 1520 279
rect 1513 272 1515 274
rect 1517 272 1520 274
rect 1513 270 1520 272
rect 1522 296 1530 298
rect 1522 294 1525 296
rect 1527 294 1530 296
rect 1522 289 1530 294
rect 1522 287 1525 289
rect 1527 287 1530 289
rect 1522 270 1530 287
rect 1532 288 1540 298
rect 1532 286 1535 288
rect 1537 286 1540 288
rect 1532 281 1540 286
rect 1532 279 1535 281
rect 1537 279 1540 281
rect 1532 270 1540 279
rect 1542 296 1556 298
rect 1542 294 1547 296
rect 1549 295 1556 296
rect 1579 296 1588 298
rect 1549 294 1558 295
rect 1542 289 1558 294
rect 1542 287 1547 289
rect 1549 287 1558 289
rect 1542 270 1558 287
rect 1560 270 1565 295
rect 1567 286 1572 295
rect 1579 294 1582 296
rect 1584 294 1588 296
rect 1579 286 1588 294
rect 1567 277 1575 286
rect 1567 275 1570 277
rect 1572 275 1575 277
rect 1567 273 1575 275
rect 1577 273 1588 286
rect 1590 286 1595 298
rect 1604 291 1609 298
rect 1602 289 1609 291
rect 1602 287 1604 289
rect 1606 287 1609 289
rect 1590 284 1597 286
rect 1602 285 1609 287
rect 1590 282 1593 284
rect 1595 282 1597 284
rect 1590 277 1597 282
rect 1604 277 1609 285
rect 1611 277 1616 298
rect 1618 296 1627 298
rect 1618 294 1623 296
rect 1625 294 1627 296
rect 1618 288 1627 294
rect 1650 289 1657 291
rect 1618 277 1629 288
rect 1590 275 1593 277
rect 1595 275 1597 277
rect 1590 273 1597 275
rect 1567 270 1572 273
rect 1621 270 1629 277
rect 1631 286 1638 288
rect 1631 284 1634 286
rect 1636 284 1638 286
rect 1631 279 1638 284
rect 1631 277 1634 279
rect 1636 277 1638 279
rect 1650 287 1652 289
rect 1654 287 1657 289
rect 1650 278 1657 287
rect 1659 289 1667 291
rect 1659 287 1662 289
rect 1664 287 1667 289
rect 1659 282 1667 287
rect 1659 280 1662 282
rect 1664 280 1667 282
rect 1659 278 1667 280
rect 1669 289 1675 291
rect 1669 287 1677 289
rect 1669 285 1672 287
rect 1674 285 1677 287
rect 1669 278 1677 285
rect 1631 275 1638 277
rect 1631 270 1636 275
rect 1671 271 1677 278
rect 1679 284 1684 289
rect 1692 286 1697 298
rect 1690 284 1697 286
rect 1679 282 1686 284
rect 1679 280 1682 282
rect 1684 280 1686 282
rect 1679 275 1686 280
rect 1679 273 1682 275
rect 1684 273 1686 275
rect 1690 282 1692 284
rect 1694 282 1697 284
rect 1690 277 1697 282
rect 1690 275 1692 277
rect 1694 275 1697 277
rect 1690 273 1697 275
rect 1699 296 1708 298
rect 1699 294 1703 296
rect 1705 294 1708 296
rect 1731 296 1745 298
rect 1731 295 1738 296
rect 1699 286 1708 294
rect 1715 286 1720 295
rect 1699 273 1710 286
rect 1712 277 1720 286
rect 1712 275 1715 277
rect 1717 275 1720 277
rect 1712 273 1720 275
rect 1679 271 1686 273
rect 1715 270 1720 273
rect 1722 270 1727 295
rect 1729 294 1738 295
rect 1740 294 1745 296
rect 1729 289 1745 294
rect 1729 287 1738 289
rect 1740 287 1745 289
rect 1729 270 1745 287
rect 1747 288 1755 298
rect 1747 286 1750 288
rect 1752 286 1755 288
rect 1747 281 1755 286
rect 1747 279 1750 281
rect 1752 279 1755 281
rect 1747 270 1755 279
rect 1757 296 1765 298
rect 1757 294 1760 296
rect 1762 294 1765 296
rect 1757 289 1765 294
rect 1757 287 1760 289
rect 1762 287 1765 289
rect 1757 270 1765 287
rect 1767 283 1772 298
rect 1782 283 1787 298
rect 1767 281 1774 283
rect 1767 279 1770 281
rect 1772 279 1774 281
rect 1767 274 1774 279
rect 1767 272 1770 274
rect 1772 272 1774 274
rect 1767 270 1774 272
rect 1780 281 1787 283
rect 1780 279 1782 281
rect 1784 279 1787 281
rect 1780 274 1787 279
rect 1780 272 1782 274
rect 1784 272 1787 274
rect 1780 270 1787 272
rect 1789 296 1797 298
rect 1789 294 1792 296
rect 1794 294 1797 296
rect 1789 289 1797 294
rect 1789 287 1792 289
rect 1794 287 1797 289
rect 1789 270 1797 287
rect 1799 288 1807 298
rect 1799 286 1802 288
rect 1804 286 1807 288
rect 1799 281 1807 286
rect 1799 279 1802 281
rect 1804 279 1807 281
rect 1799 270 1807 279
rect 1809 296 1823 298
rect 1809 294 1814 296
rect 1816 295 1823 296
rect 1846 296 1855 298
rect 1816 294 1825 295
rect 1809 289 1825 294
rect 1809 287 1814 289
rect 1816 287 1825 289
rect 1809 270 1825 287
rect 1827 270 1832 295
rect 1834 286 1839 295
rect 1846 294 1849 296
rect 1851 294 1855 296
rect 1846 286 1855 294
rect 1834 277 1842 286
rect 1834 275 1837 277
rect 1839 275 1842 277
rect 1834 273 1842 275
rect 1844 273 1855 286
rect 1857 286 1862 298
rect 1871 291 1876 298
rect 1869 289 1876 291
rect 1869 287 1871 289
rect 1873 287 1876 289
rect 1857 284 1864 286
rect 1869 285 1876 287
rect 1857 282 1860 284
rect 1862 282 1864 284
rect 1857 277 1864 282
rect 1871 277 1876 285
rect 1878 277 1883 298
rect 1885 296 1894 298
rect 1885 294 1890 296
rect 1892 294 1894 296
rect 1885 288 1894 294
rect 1885 277 1896 288
rect 1857 275 1860 277
rect 1862 275 1864 277
rect 1857 273 1864 275
rect 1834 270 1839 273
rect 1888 270 1896 277
rect 1898 286 1905 288
rect 1898 284 1901 286
rect 1903 284 1905 286
rect 1898 279 1905 284
rect 1898 277 1901 279
rect 1903 277 1905 279
rect 1922 277 1927 298
rect 1898 275 1905 277
rect 1920 275 1927 277
rect 1898 270 1903 275
rect 1920 273 1922 275
rect 1924 273 1927 275
rect 1920 271 1927 273
rect 1929 296 1941 298
rect 1929 294 1932 296
rect 1934 294 1941 296
rect 1929 289 1941 294
rect 1958 289 1963 298
rect 1929 287 1932 289
rect 1934 287 1943 289
rect 1929 271 1943 287
rect 1945 282 1953 289
rect 1945 280 1948 282
rect 1950 280 1953 282
rect 1945 275 1953 280
rect 1945 273 1948 275
rect 1950 273 1953 275
rect 1945 271 1953 273
rect 1955 282 1963 289
rect 1955 280 1958 282
rect 1960 280 1963 282
rect 1955 271 1963 280
rect 1965 292 1970 298
rect 1965 290 1972 292
rect 1965 288 1968 290
rect 1970 288 1972 290
rect 1965 286 1972 288
rect 1978 286 1983 298
rect 1965 271 1970 286
rect 1976 284 1983 286
rect 1976 282 1978 284
rect 1980 282 1983 284
rect 1976 277 1983 282
rect 1976 275 1978 277
rect 1980 275 1983 277
rect 1976 273 1983 275
rect 1985 296 1994 298
rect 1985 294 1989 296
rect 1991 294 1994 296
rect 2017 296 2031 298
rect 2017 295 2024 296
rect 1985 286 1994 294
rect 2001 286 2006 295
rect 1985 273 1996 286
rect 1998 277 2006 286
rect 1998 275 2001 277
rect 2003 275 2006 277
rect 1998 273 2006 275
rect 2001 270 2006 273
rect 2008 270 2013 295
rect 2015 294 2024 295
rect 2026 294 2031 296
rect 2015 289 2031 294
rect 2015 287 2024 289
rect 2026 287 2031 289
rect 2015 270 2031 287
rect 2033 288 2041 298
rect 2033 286 2036 288
rect 2038 286 2041 288
rect 2033 281 2041 286
rect 2033 279 2036 281
rect 2038 279 2041 281
rect 2033 270 2041 279
rect 2043 296 2051 298
rect 2043 294 2046 296
rect 2048 294 2051 296
rect 2043 289 2051 294
rect 2043 287 2046 289
rect 2048 287 2051 289
rect 2043 270 2051 287
rect 2053 283 2058 298
rect 2068 283 2073 298
rect 2053 281 2060 283
rect 2053 279 2056 281
rect 2058 279 2060 281
rect 2053 274 2060 279
rect 2053 272 2056 274
rect 2058 272 2060 274
rect 2053 270 2060 272
rect 2066 281 2073 283
rect 2066 279 2068 281
rect 2070 279 2073 281
rect 2066 274 2073 279
rect 2066 272 2068 274
rect 2070 272 2073 274
rect 2066 270 2073 272
rect 2075 296 2083 298
rect 2075 294 2078 296
rect 2080 294 2083 296
rect 2075 289 2083 294
rect 2075 287 2078 289
rect 2080 287 2083 289
rect 2075 270 2083 287
rect 2085 288 2093 298
rect 2085 286 2088 288
rect 2090 286 2093 288
rect 2085 281 2093 286
rect 2085 279 2088 281
rect 2090 279 2093 281
rect 2085 270 2093 279
rect 2095 296 2109 298
rect 2095 294 2100 296
rect 2102 295 2109 296
rect 2132 296 2141 298
rect 2102 294 2111 295
rect 2095 289 2111 294
rect 2095 287 2100 289
rect 2102 287 2111 289
rect 2095 270 2111 287
rect 2113 270 2118 295
rect 2120 286 2125 295
rect 2132 294 2135 296
rect 2137 294 2141 296
rect 2132 286 2141 294
rect 2120 277 2128 286
rect 2120 275 2123 277
rect 2125 275 2128 277
rect 2120 273 2128 275
rect 2130 273 2141 286
rect 2143 286 2148 298
rect 2157 291 2162 298
rect 2155 289 2162 291
rect 2155 287 2157 289
rect 2159 287 2162 289
rect 2143 284 2150 286
rect 2155 285 2162 287
rect 2143 282 2146 284
rect 2148 282 2150 284
rect 2143 277 2150 282
rect 2157 277 2162 285
rect 2164 277 2169 298
rect 2171 296 2180 298
rect 2171 294 2176 296
rect 2178 294 2180 296
rect 2209 296 2216 298
rect 2171 288 2180 294
rect 2209 294 2211 296
rect 2213 294 2216 296
rect 2171 277 2182 288
rect 2143 275 2146 277
rect 2148 275 2150 277
rect 2143 273 2150 275
rect 2120 270 2125 273
rect 2174 270 2182 277
rect 2184 286 2191 288
rect 2184 284 2187 286
rect 2189 284 2191 286
rect 2184 279 2191 284
rect 2209 286 2216 294
rect 2184 277 2187 279
rect 2189 277 2191 279
rect 2210 282 2216 286
rect 2218 282 2223 298
rect 2225 286 2233 298
rect 2225 284 2228 286
rect 2230 284 2233 286
rect 2225 282 2233 284
rect 2235 282 2240 298
rect 2242 296 2250 298
rect 2242 294 2245 296
rect 2247 294 2250 296
rect 2242 282 2250 294
rect 2210 278 2214 282
rect 2184 275 2191 277
rect 2201 276 2206 278
rect 2184 270 2189 275
rect 2199 274 2206 276
rect 2199 272 2201 274
rect 2203 272 2206 274
rect 2199 270 2206 272
rect 2208 270 2214 278
rect 2245 280 2250 282
rect 2252 291 2257 298
rect 2277 296 2284 298
rect 2277 294 2279 296
rect 2281 294 2284 296
rect 2252 289 2259 291
rect 2252 287 2255 289
rect 2257 287 2259 289
rect 2252 285 2259 287
rect 2277 286 2284 294
rect 2252 280 2257 285
rect 2278 282 2284 286
rect 2286 282 2291 298
rect 2293 286 2301 298
rect 2293 284 2296 286
rect 2298 284 2301 286
rect 2293 282 2301 284
rect 2303 282 2308 298
rect 2310 296 2318 298
rect 2310 294 2313 296
rect 2315 294 2318 296
rect 2310 282 2318 294
rect 2278 278 2282 282
rect 2269 276 2274 278
rect 2267 274 2274 276
rect 2267 272 2269 274
rect 2271 272 2274 274
rect 2267 270 2274 272
rect 2276 270 2282 278
rect 2313 280 2318 282
rect 2320 291 2325 298
rect 2320 289 2327 291
rect 2320 287 2323 289
rect 2325 287 2327 289
rect 2320 285 2327 287
rect 2320 280 2325 285
rect 29 186 35 193
rect 8 177 15 186
rect 8 175 10 177
rect 12 175 15 177
rect 8 173 15 175
rect 17 184 25 186
rect 17 182 20 184
rect 22 182 25 184
rect 17 177 25 182
rect 17 175 20 177
rect 22 175 25 177
rect 17 173 25 175
rect 27 179 35 186
rect 27 177 30 179
rect 32 177 35 179
rect 27 175 35 177
rect 37 190 44 193
rect 37 188 40 190
rect 42 188 44 190
rect 37 182 44 188
rect 69 186 75 193
rect 37 180 40 182
rect 42 180 44 182
rect 37 178 44 180
rect 37 175 42 178
rect 48 177 55 186
rect 48 175 50 177
rect 52 175 55 177
rect 27 173 33 175
rect 48 173 55 175
rect 57 184 65 186
rect 57 182 60 184
rect 62 182 65 184
rect 57 177 65 182
rect 57 175 60 177
rect 62 175 65 177
rect 57 173 65 175
rect 67 179 75 186
rect 67 177 70 179
rect 72 177 75 179
rect 67 175 75 177
rect 77 191 84 193
rect 113 191 118 194
rect 77 189 80 191
rect 82 189 84 191
rect 77 184 84 189
rect 77 182 80 184
rect 82 182 84 184
rect 77 180 84 182
rect 88 189 95 191
rect 88 187 90 189
rect 92 187 95 189
rect 88 182 95 187
rect 88 180 90 182
rect 92 180 95 182
rect 77 175 82 180
rect 88 178 95 180
rect 67 173 73 175
rect 90 166 95 178
rect 97 178 108 191
rect 110 189 118 191
rect 110 187 113 189
rect 115 187 118 189
rect 110 178 118 187
rect 97 170 106 178
rect 97 168 101 170
rect 103 168 106 170
rect 113 169 118 178
rect 120 169 125 194
rect 127 177 143 194
rect 127 175 136 177
rect 138 175 143 177
rect 127 170 143 175
rect 127 169 136 170
rect 97 166 106 168
rect 129 168 136 169
rect 138 168 143 170
rect 129 166 143 168
rect 145 185 153 194
rect 145 183 148 185
rect 150 183 153 185
rect 145 178 153 183
rect 145 176 148 178
rect 150 176 153 178
rect 145 166 153 176
rect 155 177 163 194
rect 155 175 158 177
rect 160 175 163 177
rect 155 170 163 175
rect 155 168 158 170
rect 160 168 163 170
rect 155 166 163 168
rect 165 192 172 194
rect 165 190 168 192
rect 170 190 172 192
rect 165 185 172 190
rect 165 183 168 185
rect 170 183 172 185
rect 165 181 172 183
rect 178 192 185 194
rect 178 190 180 192
rect 182 190 185 192
rect 178 185 185 190
rect 178 183 180 185
rect 182 183 185 185
rect 178 181 185 183
rect 165 166 170 181
rect 180 166 185 181
rect 187 177 195 194
rect 187 175 190 177
rect 192 175 195 177
rect 187 170 195 175
rect 187 168 190 170
rect 192 168 195 170
rect 187 166 195 168
rect 197 185 205 194
rect 197 183 200 185
rect 202 183 205 185
rect 197 178 205 183
rect 197 176 200 178
rect 202 176 205 178
rect 197 166 205 176
rect 207 177 223 194
rect 207 175 212 177
rect 214 175 223 177
rect 207 170 223 175
rect 207 168 212 170
rect 214 169 223 170
rect 225 169 230 194
rect 232 191 237 194
rect 232 189 240 191
rect 232 187 235 189
rect 237 187 240 189
rect 232 178 240 187
rect 242 178 253 191
rect 232 169 237 178
rect 244 170 253 178
rect 214 168 221 169
rect 207 166 221 168
rect 244 168 247 170
rect 249 168 253 170
rect 244 166 253 168
rect 255 189 262 191
rect 255 187 258 189
rect 260 187 262 189
rect 286 187 294 194
rect 255 182 262 187
rect 255 180 258 182
rect 260 180 262 182
rect 255 178 262 180
rect 269 179 274 187
rect 255 166 260 178
rect 267 177 274 179
rect 267 175 269 177
rect 271 175 274 177
rect 267 173 274 175
rect 269 166 274 173
rect 276 166 281 187
rect 283 176 294 187
rect 296 189 301 194
rect 296 187 303 189
rect 296 185 299 187
rect 301 185 303 187
rect 336 186 342 193
rect 296 180 303 185
rect 296 178 299 180
rect 301 178 303 180
rect 296 176 303 178
rect 315 177 322 186
rect 283 170 292 176
rect 315 175 317 177
rect 319 175 322 177
rect 315 173 322 175
rect 324 184 332 186
rect 324 182 327 184
rect 329 182 332 184
rect 324 177 332 182
rect 324 175 327 177
rect 329 175 332 177
rect 324 173 332 175
rect 334 179 342 186
rect 334 177 337 179
rect 339 177 342 179
rect 334 175 342 177
rect 344 191 351 193
rect 380 191 385 194
rect 344 189 347 191
rect 349 189 351 191
rect 344 184 351 189
rect 344 182 347 184
rect 349 182 351 184
rect 344 180 351 182
rect 355 189 362 191
rect 355 187 357 189
rect 359 187 362 189
rect 355 182 362 187
rect 355 180 357 182
rect 359 180 362 182
rect 344 175 349 180
rect 355 178 362 180
rect 334 173 340 175
rect 283 168 288 170
rect 290 168 292 170
rect 283 166 292 168
rect 357 166 362 178
rect 364 178 375 191
rect 377 189 385 191
rect 377 187 380 189
rect 382 187 385 189
rect 377 178 385 187
rect 364 170 373 178
rect 364 168 368 170
rect 370 168 373 170
rect 380 169 385 178
rect 387 169 392 194
rect 394 177 410 194
rect 394 175 403 177
rect 405 175 410 177
rect 394 170 410 175
rect 394 169 403 170
rect 364 166 373 168
rect 396 168 403 169
rect 405 168 410 170
rect 396 166 410 168
rect 412 185 420 194
rect 412 183 415 185
rect 417 183 420 185
rect 412 178 420 183
rect 412 176 415 178
rect 417 176 420 178
rect 412 166 420 176
rect 422 177 430 194
rect 422 175 425 177
rect 427 175 430 177
rect 422 170 430 175
rect 422 168 425 170
rect 427 168 430 170
rect 422 166 430 168
rect 432 192 439 194
rect 432 190 435 192
rect 437 190 439 192
rect 432 185 439 190
rect 432 183 435 185
rect 437 183 439 185
rect 432 181 439 183
rect 445 192 452 194
rect 445 190 447 192
rect 449 190 452 192
rect 445 185 452 190
rect 445 183 447 185
rect 449 183 452 185
rect 445 181 452 183
rect 432 166 437 181
rect 447 166 452 181
rect 454 177 462 194
rect 454 175 457 177
rect 459 175 462 177
rect 454 170 462 175
rect 454 168 457 170
rect 459 168 462 170
rect 454 166 462 168
rect 464 185 472 194
rect 464 183 467 185
rect 469 183 472 185
rect 464 178 472 183
rect 464 176 467 178
rect 469 176 472 178
rect 464 166 472 176
rect 474 177 490 194
rect 474 175 479 177
rect 481 175 490 177
rect 474 170 490 175
rect 474 168 479 170
rect 481 169 490 170
rect 492 169 497 194
rect 499 191 504 194
rect 499 189 507 191
rect 499 187 502 189
rect 504 187 507 189
rect 499 178 507 187
rect 509 178 520 191
rect 499 169 504 178
rect 511 170 520 178
rect 481 168 488 169
rect 474 166 488 168
rect 511 168 514 170
rect 516 168 520 170
rect 511 166 520 168
rect 522 189 529 191
rect 522 187 525 189
rect 527 187 529 189
rect 553 187 561 194
rect 522 182 529 187
rect 522 180 525 182
rect 527 180 529 182
rect 522 178 529 180
rect 536 179 541 187
rect 522 166 527 178
rect 534 177 541 179
rect 534 175 536 177
rect 538 175 541 177
rect 534 173 541 175
rect 536 166 541 173
rect 543 166 548 187
rect 550 176 561 187
rect 563 189 568 194
rect 563 187 570 189
rect 563 185 566 187
rect 568 185 570 187
rect 603 186 609 193
rect 563 180 570 185
rect 563 178 566 180
rect 568 178 570 180
rect 563 176 570 178
rect 582 177 589 186
rect 550 170 559 176
rect 582 175 584 177
rect 586 175 589 177
rect 582 173 589 175
rect 591 184 599 186
rect 591 182 594 184
rect 596 182 599 184
rect 591 177 599 182
rect 591 175 594 177
rect 596 175 599 177
rect 591 173 599 175
rect 601 179 609 186
rect 601 177 604 179
rect 606 177 609 179
rect 601 175 609 177
rect 611 191 618 193
rect 647 191 652 194
rect 611 189 614 191
rect 616 189 618 191
rect 611 184 618 189
rect 611 182 614 184
rect 616 182 618 184
rect 611 180 618 182
rect 622 189 629 191
rect 622 187 624 189
rect 626 187 629 189
rect 622 182 629 187
rect 622 180 624 182
rect 626 180 629 182
rect 611 175 616 180
rect 622 178 629 180
rect 601 173 607 175
rect 550 168 555 170
rect 557 168 559 170
rect 550 166 559 168
rect 624 166 629 178
rect 631 178 642 191
rect 644 189 652 191
rect 644 187 647 189
rect 649 187 652 189
rect 644 178 652 187
rect 631 170 640 178
rect 631 168 635 170
rect 637 168 640 170
rect 647 169 652 178
rect 654 169 659 194
rect 661 177 677 194
rect 661 175 670 177
rect 672 175 677 177
rect 661 170 677 175
rect 661 169 670 170
rect 631 166 640 168
rect 663 168 670 169
rect 672 168 677 170
rect 663 166 677 168
rect 679 185 687 194
rect 679 183 682 185
rect 684 183 687 185
rect 679 178 687 183
rect 679 176 682 178
rect 684 176 687 178
rect 679 166 687 176
rect 689 177 697 194
rect 689 175 692 177
rect 694 175 697 177
rect 689 170 697 175
rect 689 168 692 170
rect 694 168 697 170
rect 689 166 697 168
rect 699 192 706 194
rect 699 190 702 192
rect 704 190 706 192
rect 699 185 706 190
rect 699 183 702 185
rect 704 183 706 185
rect 699 181 706 183
rect 712 192 719 194
rect 712 190 714 192
rect 716 190 719 192
rect 712 185 719 190
rect 712 183 714 185
rect 716 183 719 185
rect 712 181 719 183
rect 699 166 704 181
rect 714 166 719 181
rect 721 177 729 194
rect 721 175 724 177
rect 726 175 729 177
rect 721 170 729 175
rect 721 168 724 170
rect 726 168 729 170
rect 721 166 729 168
rect 731 185 739 194
rect 731 183 734 185
rect 736 183 739 185
rect 731 178 739 183
rect 731 176 734 178
rect 736 176 739 178
rect 731 166 739 176
rect 741 177 757 194
rect 741 175 746 177
rect 748 175 757 177
rect 741 170 757 175
rect 741 168 746 170
rect 748 169 757 170
rect 759 169 764 194
rect 766 191 771 194
rect 766 189 774 191
rect 766 187 769 189
rect 771 187 774 189
rect 766 178 774 187
rect 776 178 787 191
rect 766 169 771 178
rect 778 170 787 178
rect 748 168 755 169
rect 741 166 755 168
rect 778 168 781 170
rect 783 168 787 170
rect 778 166 787 168
rect 789 189 796 191
rect 789 187 792 189
rect 794 187 796 189
rect 820 187 828 194
rect 789 182 796 187
rect 789 180 792 182
rect 794 180 796 182
rect 789 178 796 180
rect 803 179 808 187
rect 789 166 794 178
rect 801 177 808 179
rect 801 175 803 177
rect 805 175 808 177
rect 801 173 808 175
rect 803 166 808 173
rect 810 166 815 187
rect 817 176 828 187
rect 830 189 835 194
rect 830 187 837 189
rect 830 185 833 187
rect 835 185 837 187
rect 870 186 876 193
rect 830 180 837 185
rect 830 178 833 180
rect 835 178 837 180
rect 830 176 837 178
rect 849 177 856 186
rect 817 170 826 176
rect 849 175 851 177
rect 853 175 856 177
rect 849 173 856 175
rect 858 184 866 186
rect 858 182 861 184
rect 863 182 866 184
rect 858 177 866 182
rect 858 175 861 177
rect 863 175 866 177
rect 858 173 866 175
rect 868 179 876 186
rect 868 177 871 179
rect 873 177 876 179
rect 868 175 876 177
rect 878 191 885 193
rect 914 191 919 194
rect 878 189 881 191
rect 883 189 885 191
rect 878 184 885 189
rect 878 182 881 184
rect 883 182 885 184
rect 878 180 885 182
rect 889 189 896 191
rect 889 187 891 189
rect 893 187 896 189
rect 889 182 896 187
rect 889 180 891 182
rect 893 180 896 182
rect 878 175 883 180
rect 889 178 896 180
rect 868 173 874 175
rect 817 168 822 170
rect 824 168 826 170
rect 817 166 826 168
rect 891 166 896 178
rect 898 178 909 191
rect 911 189 919 191
rect 911 187 914 189
rect 916 187 919 189
rect 911 178 919 187
rect 898 170 907 178
rect 898 168 902 170
rect 904 168 907 170
rect 914 169 919 178
rect 921 169 926 194
rect 928 177 944 194
rect 928 175 937 177
rect 939 175 944 177
rect 928 170 944 175
rect 928 169 937 170
rect 898 166 907 168
rect 930 168 937 169
rect 939 168 944 170
rect 930 166 944 168
rect 946 185 954 194
rect 946 183 949 185
rect 951 183 954 185
rect 946 178 954 183
rect 946 176 949 178
rect 951 176 954 178
rect 946 166 954 176
rect 956 177 964 194
rect 956 175 959 177
rect 961 175 964 177
rect 956 170 964 175
rect 956 168 959 170
rect 961 168 964 170
rect 956 166 964 168
rect 966 192 973 194
rect 966 190 969 192
rect 971 190 973 192
rect 966 185 973 190
rect 966 183 969 185
rect 971 183 973 185
rect 966 181 973 183
rect 979 192 986 194
rect 979 190 981 192
rect 983 190 986 192
rect 979 185 986 190
rect 979 183 981 185
rect 983 183 986 185
rect 979 181 986 183
rect 966 166 971 181
rect 981 166 986 181
rect 988 177 996 194
rect 988 175 991 177
rect 993 175 996 177
rect 988 170 996 175
rect 988 168 991 170
rect 993 168 996 170
rect 988 166 996 168
rect 998 185 1006 194
rect 998 183 1001 185
rect 1003 183 1006 185
rect 998 178 1006 183
rect 998 176 1001 178
rect 1003 176 1006 178
rect 998 166 1006 176
rect 1008 177 1024 194
rect 1008 175 1013 177
rect 1015 175 1024 177
rect 1008 170 1024 175
rect 1008 168 1013 170
rect 1015 169 1024 170
rect 1026 169 1031 194
rect 1033 191 1038 194
rect 1033 189 1041 191
rect 1033 187 1036 189
rect 1038 187 1041 189
rect 1033 178 1041 187
rect 1043 178 1054 191
rect 1033 169 1038 178
rect 1045 170 1054 178
rect 1015 168 1022 169
rect 1008 166 1022 168
rect 1045 168 1048 170
rect 1050 168 1054 170
rect 1045 166 1054 168
rect 1056 189 1063 191
rect 1056 187 1059 189
rect 1061 187 1063 189
rect 1087 187 1095 194
rect 1056 182 1063 187
rect 1056 180 1059 182
rect 1061 180 1063 182
rect 1056 178 1063 180
rect 1070 179 1075 187
rect 1056 166 1061 178
rect 1068 177 1075 179
rect 1068 175 1070 177
rect 1072 175 1075 177
rect 1068 173 1075 175
rect 1070 166 1075 173
rect 1077 166 1082 187
rect 1084 176 1095 187
rect 1097 189 1102 194
rect 1097 187 1104 189
rect 1097 185 1100 187
rect 1102 185 1104 187
rect 1137 186 1143 193
rect 1097 180 1104 185
rect 1097 178 1100 180
rect 1102 178 1104 180
rect 1097 176 1104 178
rect 1116 177 1123 186
rect 1084 170 1093 176
rect 1116 175 1118 177
rect 1120 175 1123 177
rect 1116 173 1123 175
rect 1125 184 1133 186
rect 1125 182 1128 184
rect 1130 182 1133 184
rect 1125 177 1133 182
rect 1125 175 1128 177
rect 1130 175 1133 177
rect 1125 173 1133 175
rect 1135 179 1143 186
rect 1135 177 1138 179
rect 1140 177 1143 179
rect 1135 175 1143 177
rect 1145 191 1152 193
rect 1181 191 1186 194
rect 1145 189 1148 191
rect 1150 189 1152 191
rect 1145 184 1152 189
rect 1145 182 1148 184
rect 1150 182 1152 184
rect 1145 180 1152 182
rect 1156 189 1163 191
rect 1156 187 1158 189
rect 1160 187 1163 189
rect 1156 182 1163 187
rect 1156 180 1158 182
rect 1160 180 1163 182
rect 1145 175 1150 180
rect 1156 178 1163 180
rect 1135 173 1141 175
rect 1084 168 1089 170
rect 1091 168 1093 170
rect 1084 166 1093 168
rect 1158 166 1163 178
rect 1165 178 1176 191
rect 1178 189 1186 191
rect 1178 187 1181 189
rect 1183 187 1186 189
rect 1178 178 1186 187
rect 1165 170 1174 178
rect 1165 168 1169 170
rect 1171 168 1174 170
rect 1181 169 1186 178
rect 1188 169 1193 194
rect 1195 177 1211 194
rect 1195 175 1204 177
rect 1206 175 1211 177
rect 1195 170 1211 175
rect 1195 169 1204 170
rect 1165 166 1174 168
rect 1197 168 1204 169
rect 1206 168 1211 170
rect 1197 166 1211 168
rect 1213 185 1221 194
rect 1213 183 1216 185
rect 1218 183 1221 185
rect 1213 178 1221 183
rect 1213 176 1216 178
rect 1218 176 1221 178
rect 1213 166 1221 176
rect 1223 177 1231 194
rect 1223 175 1226 177
rect 1228 175 1231 177
rect 1223 170 1231 175
rect 1223 168 1226 170
rect 1228 168 1231 170
rect 1223 166 1231 168
rect 1233 192 1240 194
rect 1233 190 1236 192
rect 1238 190 1240 192
rect 1233 185 1240 190
rect 1233 183 1236 185
rect 1238 183 1240 185
rect 1233 181 1240 183
rect 1246 192 1253 194
rect 1246 190 1248 192
rect 1250 190 1253 192
rect 1246 185 1253 190
rect 1246 183 1248 185
rect 1250 183 1253 185
rect 1246 181 1253 183
rect 1233 166 1238 181
rect 1248 166 1253 181
rect 1255 177 1263 194
rect 1255 175 1258 177
rect 1260 175 1263 177
rect 1255 170 1263 175
rect 1255 168 1258 170
rect 1260 168 1263 170
rect 1255 166 1263 168
rect 1265 185 1273 194
rect 1265 183 1268 185
rect 1270 183 1273 185
rect 1265 178 1273 183
rect 1265 176 1268 178
rect 1270 176 1273 178
rect 1265 166 1273 176
rect 1275 177 1291 194
rect 1275 175 1280 177
rect 1282 175 1291 177
rect 1275 170 1291 175
rect 1275 168 1280 170
rect 1282 169 1291 170
rect 1293 169 1298 194
rect 1300 191 1305 194
rect 1300 189 1308 191
rect 1300 187 1303 189
rect 1305 187 1308 189
rect 1300 178 1308 187
rect 1310 178 1321 191
rect 1300 169 1305 178
rect 1312 170 1321 178
rect 1282 168 1289 169
rect 1275 166 1289 168
rect 1312 168 1315 170
rect 1317 168 1321 170
rect 1312 166 1321 168
rect 1323 189 1330 191
rect 1323 187 1326 189
rect 1328 187 1330 189
rect 1354 187 1362 194
rect 1323 182 1330 187
rect 1323 180 1326 182
rect 1328 180 1330 182
rect 1323 178 1330 180
rect 1337 179 1342 187
rect 1323 166 1328 178
rect 1335 177 1342 179
rect 1335 175 1337 177
rect 1339 175 1342 177
rect 1335 173 1342 175
rect 1337 166 1342 173
rect 1344 166 1349 187
rect 1351 176 1362 187
rect 1364 189 1369 194
rect 1364 187 1371 189
rect 1364 185 1367 187
rect 1369 185 1371 187
rect 1404 186 1410 193
rect 1364 180 1371 185
rect 1364 178 1367 180
rect 1369 178 1371 180
rect 1364 176 1371 178
rect 1383 177 1390 186
rect 1351 170 1360 176
rect 1383 175 1385 177
rect 1387 175 1390 177
rect 1383 173 1390 175
rect 1392 184 1400 186
rect 1392 182 1395 184
rect 1397 182 1400 184
rect 1392 177 1400 182
rect 1392 175 1395 177
rect 1397 175 1400 177
rect 1392 173 1400 175
rect 1402 179 1410 186
rect 1402 177 1405 179
rect 1407 177 1410 179
rect 1402 175 1410 177
rect 1412 191 1419 193
rect 1448 191 1453 194
rect 1412 189 1415 191
rect 1417 189 1419 191
rect 1412 184 1419 189
rect 1412 182 1415 184
rect 1417 182 1419 184
rect 1412 180 1419 182
rect 1423 189 1430 191
rect 1423 187 1425 189
rect 1427 187 1430 189
rect 1423 182 1430 187
rect 1423 180 1425 182
rect 1427 180 1430 182
rect 1412 175 1417 180
rect 1423 178 1430 180
rect 1402 173 1408 175
rect 1351 168 1356 170
rect 1358 168 1360 170
rect 1351 166 1360 168
rect 1425 166 1430 178
rect 1432 178 1443 191
rect 1445 189 1453 191
rect 1445 187 1448 189
rect 1450 187 1453 189
rect 1445 178 1453 187
rect 1432 170 1441 178
rect 1432 168 1436 170
rect 1438 168 1441 170
rect 1448 169 1453 178
rect 1455 169 1460 194
rect 1462 177 1478 194
rect 1462 175 1471 177
rect 1473 175 1478 177
rect 1462 170 1478 175
rect 1462 169 1471 170
rect 1432 166 1441 168
rect 1464 168 1471 169
rect 1473 168 1478 170
rect 1464 166 1478 168
rect 1480 185 1488 194
rect 1480 183 1483 185
rect 1485 183 1488 185
rect 1480 178 1488 183
rect 1480 176 1483 178
rect 1485 176 1488 178
rect 1480 166 1488 176
rect 1490 177 1498 194
rect 1490 175 1493 177
rect 1495 175 1498 177
rect 1490 170 1498 175
rect 1490 168 1493 170
rect 1495 168 1498 170
rect 1490 166 1498 168
rect 1500 192 1507 194
rect 1500 190 1503 192
rect 1505 190 1507 192
rect 1500 185 1507 190
rect 1500 183 1503 185
rect 1505 183 1507 185
rect 1500 181 1507 183
rect 1513 192 1520 194
rect 1513 190 1515 192
rect 1517 190 1520 192
rect 1513 185 1520 190
rect 1513 183 1515 185
rect 1517 183 1520 185
rect 1513 181 1520 183
rect 1500 166 1505 181
rect 1515 166 1520 181
rect 1522 177 1530 194
rect 1522 175 1525 177
rect 1527 175 1530 177
rect 1522 170 1530 175
rect 1522 168 1525 170
rect 1527 168 1530 170
rect 1522 166 1530 168
rect 1532 185 1540 194
rect 1532 183 1535 185
rect 1537 183 1540 185
rect 1532 178 1540 183
rect 1532 176 1535 178
rect 1537 176 1540 178
rect 1532 166 1540 176
rect 1542 177 1558 194
rect 1542 175 1547 177
rect 1549 175 1558 177
rect 1542 170 1558 175
rect 1542 168 1547 170
rect 1549 169 1558 170
rect 1560 169 1565 194
rect 1567 191 1572 194
rect 1567 189 1575 191
rect 1567 187 1570 189
rect 1572 187 1575 189
rect 1567 178 1575 187
rect 1577 178 1588 191
rect 1567 169 1572 178
rect 1579 170 1588 178
rect 1549 168 1556 169
rect 1542 166 1556 168
rect 1579 168 1582 170
rect 1584 168 1588 170
rect 1579 166 1588 168
rect 1590 189 1597 191
rect 1590 187 1593 189
rect 1595 187 1597 189
rect 1621 187 1629 194
rect 1590 182 1597 187
rect 1590 180 1593 182
rect 1595 180 1597 182
rect 1590 178 1597 180
rect 1604 179 1609 187
rect 1590 166 1595 178
rect 1602 177 1609 179
rect 1602 175 1604 177
rect 1606 175 1609 177
rect 1602 173 1609 175
rect 1604 166 1609 173
rect 1611 166 1616 187
rect 1618 176 1629 187
rect 1631 189 1636 194
rect 1631 187 1638 189
rect 1631 185 1634 187
rect 1636 185 1638 187
rect 1671 186 1677 193
rect 1631 180 1638 185
rect 1631 178 1634 180
rect 1636 178 1638 180
rect 1631 176 1638 178
rect 1650 177 1657 186
rect 1618 170 1627 176
rect 1650 175 1652 177
rect 1654 175 1657 177
rect 1650 173 1657 175
rect 1659 184 1667 186
rect 1659 182 1662 184
rect 1664 182 1667 184
rect 1659 177 1667 182
rect 1659 175 1662 177
rect 1664 175 1667 177
rect 1659 173 1667 175
rect 1669 179 1677 186
rect 1669 177 1672 179
rect 1674 177 1677 179
rect 1669 175 1677 177
rect 1679 191 1686 193
rect 1715 191 1720 194
rect 1679 189 1682 191
rect 1684 189 1686 191
rect 1679 184 1686 189
rect 1679 182 1682 184
rect 1684 182 1686 184
rect 1679 180 1686 182
rect 1690 189 1697 191
rect 1690 187 1692 189
rect 1694 187 1697 189
rect 1690 182 1697 187
rect 1690 180 1692 182
rect 1694 180 1697 182
rect 1679 175 1684 180
rect 1690 178 1697 180
rect 1669 173 1675 175
rect 1618 168 1623 170
rect 1625 168 1627 170
rect 1618 166 1627 168
rect 1692 166 1697 178
rect 1699 178 1710 191
rect 1712 189 1720 191
rect 1712 187 1715 189
rect 1717 187 1720 189
rect 1712 178 1720 187
rect 1699 170 1708 178
rect 1699 168 1703 170
rect 1705 168 1708 170
rect 1715 169 1720 178
rect 1722 169 1727 194
rect 1729 177 1745 194
rect 1729 175 1738 177
rect 1740 175 1745 177
rect 1729 170 1745 175
rect 1729 169 1738 170
rect 1699 166 1708 168
rect 1731 168 1738 169
rect 1740 168 1745 170
rect 1731 166 1745 168
rect 1747 185 1755 194
rect 1747 183 1750 185
rect 1752 183 1755 185
rect 1747 178 1755 183
rect 1747 176 1750 178
rect 1752 176 1755 178
rect 1747 166 1755 176
rect 1757 177 1765 194
rect 1757 175 1760 177
rect 1762 175 1765 177
rect 1757 170 1765 175
rect 1757 168 1760 170
rect 1762 168 1765 170
rect 1757 166 1765 168
rect 1767 192 1774 194
rect 1767 190 1770 192
rect 1772 190 1774 192
rect 1767 185 1774 190
rect 1767 183 1770 185
rect 1772 183 1774 185
rect 1767 181 1774 183
rect 1780 192 1787 194
rect 1780 190 1782 192
rect 1784 190 1787 192
rect 1780 185 1787 190
rect 1780 183 1782 185
rect 1784 183 1787 185
rect 1780 181 1787 183
rect 1767 166 1772 181
rect 1782 166 1787 181
rect 1789 177 1797 194
rect 1789 175 1792 177
rect 1794 175 1797 177
rect 1789 170 1797 175
rect 1789 168 1792 170
rect 1794 168 1797 170
rect 1789 166 1797 168
rect 1799 185 1807 194
rect 1799 183 1802 185
rect 1804 183 1807 185
rect 1799 178 1807 183
rect 1799 176 1802 178
rect 1804 176 1807 178
rect 1799 166 1807 176
rect 1809 177 1825 194
rect 1809 175 1814 177
rect 1816 175 1825 177
rect 1809 170 1825 175
rect 1809 168 1814 170
rect 1816 169 1825 170
rect 1827 169 1832 194
rect 1834 191 1839 194
rect 1834 189 1842 191
rect 1834 187 1837 189
rect 1839 187 1842 189
rect 1834 178 1842 187
rect 1844 178 1855 191
rect 1834 169 1839 178
rect 1846 170 1855 178
rect 1816 168 1823 169
rect 1809 166 1823 168
rect 1846 168 1849 170
rect 1851 168 1855 170
rect 1846 166 1855 168
rect 1857 189 1864 191
rect 1857 187 1860 189
rect 1862 187 1864 189
rect 1888 187 1896 194
rect 1857 182 1864 187
rect 1857 180 1860 182
rect 1862 180 1864 182
rect 1857 178 1864 180
rect 1871 179 1876 187
rect 1857 166 1862 178
rect 1869 177 1876 179
rect 1869 175 1871 177
rect 1873 175 1876 177
rect 1869 173 1876 175
rect 1871 166 1876 173
rect 1878 166 1883 187
rect 1885 176 1896 187
rect 1898 189 1903 194
rect 1920 191 1927 193
rect 1920 189 1922 191
rect 1924 189 1927 191
rect 1898 187 1905 189
rect 1920 187 1927 189
rect 1898 185 1901 187
rect 1903 185 1905 187
rect 1898 180 1905 185
rect 1898 178 1901 180
rect 1903 178 1905 180
rect 1898 176 1905 178
rect 1885 170 1894 176
rect 1885 168 1890 170
rect 1892 168 1894 170
rect 1885 166 1894 168
rect 1922 166 1927 187
rect 1929 177 1943 193
rect 1929 175 1932 177
rect 1934 175 1943 177
rect 1945 191 1953 193
rect 1945 189 1948 191
rect 1950 189 1953 191
rect 1945 184 1953 189
rect 1945 182 1948 184
rect 1950 182 1953 184
rect 1945 175 1953 182
rect 1955 184 1963 193
rect 1955 182 1958 184
rect 1960 182 1963 184
rect 1955 175 1963 182
rect 1929 170 1941 175
rect 1929 168 1932 170
rect 1934 168 1941 170
rect 1929 166 1941 168
rect 1958 166 1963 175
rect 1965 178 1970 193
rect 2001 191 2006 194
rect 1976 189 1983 191
rect 1976 187 1978 189
rect 1980 187 1983 189
rect 1976 182 1983 187
rect 1976 180 1978 182
rect 1980 180 1983 182
rect 1976 178 1983 180
rect 1965 176 1972 178
rect 1965 174 1968 176
rect 1970 174 1972 176
rect 1965 172 1972 174
rect 1965 166 1970 172
rect 1978 166 1983 178
rect 1985 178 1996 191
rect 1998 189 2006 191
rect 1998 187 2001 189
rect 2003 187 2006 189
rect 1998 178 2006 187
rect 1985 170 1994 178
rect 1985 168 1989 170
rect 1991 168 1994 170
rect 2001 169 2006 178
rect 2008 169 2013 194
rect 2015 177 2031 194
rect 2015 175 2024 177
rect 2026 175 2031 177
rect 2015 170 2031 175
rect 2015 169 2024 170
rect 1985 166 1994 168
rect 2017 168 2024 169
rect 2026 168 2031 170
rect 2017 166 2031 168
rect 2033 185 2041 194
rect 2033 183 2036 185
rect 2038 183 2041 185
rect 2033 178 2041 183
rect 2033 176 2036 178
rect 2038 176 2041 178
rect 2033 166 2041 176
rect 2043 177 2051 194
rect 2043 175 2046 177
rect 2048 175 2051 177
rect 2043 170 2051 175
rect 2043 168 2046 170
rect 2048 168 2051 170
rect 2043 166 2051 168
rect 2053 192 2060 194
rect 2053 190 2056 192
rect 2058 190 2060 192
rect 2053 185 2060 190
rect 2053 183 2056 185
rect 2058 183 2060 185
rect 2053 181 2060 183
rect 2066 192 2073 194
rect 2066 190 2068 192
rect 2070 190 2073 192
rect 2066 185 2073 190
rect 2066 183 2068 185
rect 2070 183 2073 185
rect 2066 181 2073 183
rect 2053 166 2058 181
rect 2068 166 2073 181
rect 2075 177 2083 194
rect 2075 175 2078 177
rect 2080 175 2083 177
rect 2075 170 2083 175
rect 2075 168 2078 170
rect 2080 168 2083 170
rect 2075 166 2083 168
rect 2085 185 2093 194
rect 2085 183 2088 185
rect 2090 183 2093 185
rect 2085 178 2093 183
rect 2085 176 2088 178
rect 2090 176 2093 178
rect 2085 166 2093 176
rect 2095 177 2111 194
rect 2095 175 2100 177
rect 2102 175 2111 177
rect 2095 170 2111 175
rect 2095 168 2100 170
rect 2102 169 2111 170
rect 2113 169 2118 194
rect 2120 191 2125 194
rect 2120 189 2128 191
rect 2120 187 2123 189
rect 2125 187 2128 189
rect 2120 178 2128 187
rect 2130 178 2141 191
rect 2120 169 2125 178
rect 2132 170 2141 178
rect 2102 168 2109 169
rect 2095 166 2109 168
rect 2132 168 2135 170
rect 2137 168 2141 170
rect 2132 166 2141 168
rect 2143 189 2150 191
rect 2143 187 2146 189
rect 2148 187 2150 189
rect 2174 187 2182 194
rect 2143 182 2150 187
rect 2143 180 2146 182
rect 2148 180 2150 182
rect 2143 178 2150 180
rect 2157 179 2162 187
rect 2143 166 2148 178
rect 2155 177 2162 179
rect 2155 175 2157 177
rect 2159 175 2162 177
rect 2155 173 2162 175
rect 2157 166 2162 173
rect 2164 166 2169 187
rect 2171 176 2182 187
rect 2184 189 2189 194
rect 2199 192 2206 194
rect 2199 190 2201 192
rect 2203 190 2206 192
rect 2184 187 2191 189
rect 2199 188 2206 190
rect 2184 185 2187 187
rect 2189 185 2191 187
rect 2201 186 2206 188
rect 2208 186 2214 194
rect 2184 180 2191 185
rect 2184 178 2187 180
rect 2189 178 2191 180
rect 2184 176 2191 178
rect 2210 182 2214 186
rect 2267 192 2274 194
rect 2267 190 2269 192
rect 2271 190 2274 192
rect 2267 188 2274 190
rect 2269 186 2274 188
rect 2276 186 2282 194
rect 2245 182 2250 184
rect 2210 178 2216 182
rect 2171 170 2180 176
rect 2171 168 2176 170
rect 2178 168 2180 170
rect 2209 170 2216 178
rect 2171 166 2180 168
rect 2209 168 2211 170
rect 2213 168 2216 170
rect 2209 166 2216 168
rect 2218 166 2223 182
rect 2225 180 2233 182
rect 2225 178 2228 180
rect 2230 178 2233 180
rect 2225 166 2233 178
rect 2235 166 2240 182
rect 2242 170 2250 182
rect 2242 168 2245 170
rect 2247 168 2250 170
rect 2242 166 2250 168
rect 2252 179 2257 184
rect 2278 182 2282 186
rect 2313 182 2318 184
rect 2252 177 2259 179
rect 2278 178 2284 182
rect 2252 175 2255 177
rect 2257 175 2259 177
rect 2252 173 2259 175
rect 2252 166 2257 173
rect 2277 170 2284 178
rect 2277 168 2279 170
rect 2281 168 2284 170
rect 2277 166 2284 168
rect 2286 166 2291 182
rect 2293 180 2301 182
rect 2293 178 2296 180
rect 2298 178 2301 180
rect 2293 166 2301 178
rect 2303 166 2308 182
rect 2310 170 2318 182
rect 2310 168 2313 170
rect 2315 168 2318 170
rect 2310 166 2318 168
rect 2320 179 2325 184
rect 2320 177 2327 179
rect 2320 175 2323 177
rect 2325 175 2327 177
rect 2320 173 2327 175
rect 2320 166 2325 173
rect 8 145 15 147
rect 8 143 10 145
rect 12 143 15 145
rect 8 134 15 143
rect 17 145 25 147
rect 17 143 20 145
rect 22 143 25 145
rect 17 138 25 143
rect 17 136 20 138
rect 22 136 25 138
rect 17 134 25 136
rect 27 145 33 147
rect 48 145 55 147
rect 27 143 35 145
rect 27 141 30 143
rect 32 141 35 143
rect 27 134 35 141
rect 29 127 35 134
rect 37 143 42 145
rect 48 143 50 145
rect 52 143 55 145
rect 37 141 44 143
rect 37 139 40 141
rect 42 139 44 141
rect 37 133 44 139
rect 48 134 55 143
rect 57 145 65 147
rect 57 143 60 145
rect 62 143 65 145
rect 57 138 65 143
rect 57 136 60 138
rect 62 136 65 138
rect 57 134 65 136
rect 67 145 73 147
rect 67 143 75 145
rect 67 141 70 143
rect 72 141 75 143
rect 67 134 75 141
rect 37 131 40 133
rect 42 131 44 133
rect 37 127 44 131
rect 69 127 75 134
rect 77 140 82 145
rect 90 142 95 154
rect 88 140 95 142
rect 77 138 84 140
rect 77 136 80 138
rect 82 136 84 138
rect 77 131 84 136
rect 77 129 80 131
rect 82 129 84 131
rect 88 138 90 140
rect 92 138 95 140
rect 88 133 95 138
rect 88 131 90 133
rect 92 131 95 133
rect 88 129 95 131
rect 97 152 106 154
rect 97 150 101 152
rect 103 150 106 152
rect 129 152 143 154
rect 129 151 136 152
rect 97 142 106 150
rect 113 142 118 151
rect 97 129 108 142
rect 110 133 118 142
rect 110 131 113 133
rect 115 131 118 133
rect 110 129 118 131
rect 77 127 84 129
rect 113 126 118 129
rect 120 126 125 151
rect 127 150 136 151
rect 138 150 143 152
rect 127 145 143 150
rect 127 143 136 145
rect 138 143 143 145
rect 127 126 143 143
rect 145 144 153 154
rect 145 142 148 144
rect 150 142 153 144
rect 145 137 153 142
rect 145 135 148 137
rect 150 135 153 137
rect 145 126 153 135
rect 155 152 163 154
rect 155 150 158 152
rect 160 150 163 152
rect 155 145 163 150
rect 155 143 158 145
rect 160 143 163 145
rect 155 126 163 143
rect 165 139 170 154
rect 180 139 185 154
rect 165 137 172 139
rect 165 135 168 137
rect 170 135 172 137
rect 165 130 172 135
rect 165 128 168 130
rect 170 128 172 130
rect 165 126 172 128
rect 178 137 185 139
rect 178 135 180 137
rect 182 135 185 137
rect 178 130 185 135
rect 178 128 180 130
rect 182 128 185 130
rect 178 126 185 128
rect 187 152 195 154
rect 187 150 190 152
rect 192 150 195 152
rect 187 145 195 150
rect 187 143 190 145
rect 192 143 195 145
rect 187 126 195 143
rect 197 144 205 154
rect 197 142 200 144
rect 202 142 205 144
rect 197 137 205 142
rect 197 135 200 137
rect 202 135 205 137
rect 197 126 205 135
rect 207 152 221 154
rect 207 150 212 152
rect 214 151 221 152
rect 244 152 253 154
rect 214 150 223 151
rect 207 145 223 150
rect 207 143 212 145
rect 214 143 223 145
rect 207 126 223 143
rect 225 126 230 151
rect 232 142 237 151
rect 244 150 247 152
rect 249 150 253 152
rect 244 142 253 150
rect 232 133 240 142
rect 232 131 235 133
rect 237 131 240 133
rect 232 129 240 131
rect 242 129 253 142
rect 255 142 260 154
rect 269 147 274 154
rect 267 145 274 147
rect 267 143 269 145
rect 271 143 274 145
rect 255 140 262 142
rect 267 141 274 143
rect 255 138 258 140
rect 260 138 262 140
rect 255 133 262 138
rect 269 133 274 141
rect 276 133 281 154
rect 283 152 292 154
rect 283 150 288 152
rect 290 150 292 152
rect 283 144 292 150
rect 315 145 322 147
rect 283 133 294 144
rect 255 131 258 133
rect 260 131 262 133
rect 255 129 262 131
rect 232 126 237 129
rect 286 126 294 133
rect 296 142 303 144
rect 296 140 299 142
rect 301 140 303 142
rect 296 135 303 140
rect 296 133 299 135
rect 301 133 303 135
rect 315 143 317 145
rect 319 143 322 145
rect 315 134 322 143
rect 324 145 332 147
rect 324 143 327 145
rect 329 143 332 145
rect 324 138 332 143
rect 324 136 327 138
rect 329 136 332 138
rect 324 134 332 136
rect 334 145 340 147
rect 334 143 342 145
rect 334 141 337 143
rect 339 141 342 143
rect 334 134 342 141
rect 296 131 303 133
rect 296 126 301 131
rect 336 127 342 134
rect 344 140 349 145
rect 357 142 362 154
rect 355 140 362 142
rect 344 138 351 140
rect 344 136 347 138
rect 349 136 351 138
rect 344 131 351 136
rect 344 129 347 131
rect 349 129 351 131
rect 355 138 357 140
rect 359 138 362 140
rect 355 133 362 138
rect 355 131 357 133
rect 359 131 362 133
rect 355 129 362 131
rect 364 152 373 154
rect 364 150 368 152
rect 370 150 373 152
rect 396 152 410 154
rect 396 151 403 152
rect 364 142 373 150
rect 380 142 385 151
rect 364 129 375 142
rect 377 133 385 142
rect 377 131 380 133
rect 382 131 385 133
rect 377 129 385 131
rect 344 127 351 129
rect 380 126 385 129
rect 387 126 392 151
rect 394 150 403 151
rect 405 150 410 152
rect 394 145 410 150
rect 394 143 403 145
rect 405 143 410 145
rect 394 126 410 143
rect 412 144 420 154
rect 412 142 415 144
rect 417 142 420 144
rect 412 137 420 142
rect 412 135 415 137
rect 417 135 420 137
rect 412 126 420 135
rect 422 152 430 154
rect 422 150 425 152
rect 427 150 430 152
rect 422 145 430 150
rect 422 143 425 145
rect 427 143 430 145
rect 422 126 430 143
rect 432 139 437 154
rect 447 139 452 154
rect 432 137 439 139
rect 432 135 435 137
rect 437 135 439 137
rect 432 130 439 135
rect 432 128 435 130
rect 437 128 439 130
rect 432 126 439 128
rect 445 137 452 139
rect 445 135 447 137
rect 449 135 452 137
rect 445 130 452 135
rect 445 128 447 130
rect 449 128 452 130
rect 445 126 452 128
rect 454 152 462 154
rect 454 150 457 152
rect 459 150 462 152
rect 454 145 462 150
rect 454 143 457 145
rect 459 143 462 145
rect 454 126 462 143
rect 464 144 472 154
rect 464 142 467 144
rect 469 142 472 144
rect 464 137 472 142
rect 464 135 467 137
rect 469 135 472 137
rect 464 126 472 135
rect 474 152 488 154
rect 474 150 479 152
rect 481 151 488 152
rect 511 152 520 154
rect 481 150 490 151
rect 474 145 490 150
rect 474 143 479 145
rect 481 143 490 145
rect 474 126 490 143
rect 492 126 497 151
rect 499 142 504 151
rect 511 150 514 152
rect 516 150 520 152
rect 511 142 520 150
rect 499 133 507 142
rect 499 131 502 133
rect 504 131 507 133
rect 499 129 507 131
rect 509 129 520 142
rect 522 142 527 154
rect 536 147 541 154
rect 534 145 541 147
rect 534 143 536 145
rect 538 143 541 145
rect 522 140 529 142
rect 534 141 541 143
rect 522 138 525 140
rect 527 138 529 140
rect 522 133 529 138
rect 536 133 541 141
rect 543 133 548 154
rect 550 152 559 154
rect 550 150 555 152
rect 557 150 559 152
rect 550 144 559 150
rect 582 145 589 147
rect 550 133 561 144
rect 522 131 525 133
rect 527 131 529 133
rect 522 129 529 131
rect 499 126 504 129
rect 553 126 561 133
rect 563 142 570 144
rect 563 140 566 142
rect 568 140 570 142
rect 563 135 570 140
rect 563 133 566 135
rect 568 133 570 135
rect 582 143 584 145
rect 586 143 589 145
rect 582 134 589 143
rect 591 145 599 147
rect 591 143 594 145
rect 596 143 599 145
rect 591 138 599 143
rect 591 136 594 138
rect 596 136 599 138
rect 591 134 599 136
rect 601 145 607 147
rect 601 143 609 145
rect 601 141 604 143
rect 606 141 609 143
rect 601 134 609 141
rect 563 131 570 133
rect 563 126 568 131
rect 603 127 609 134
rect 611 140 616 145
rect 624 142 629 154
rect 622 140 629 142
rect 611 138 618 140
rect 611 136 614 138
rect 616 136 618 138
rect 611 131 618 136
rect 611 129 614 131
rect 616 129 618 131
rect 622 138 624 140
rect 626 138 629 140
rect 622 133 629 138
rect 622 131 624 133
rect 626 131 629 133
rect 622 129 629 131
rect 631 152 640 154
rect 631 150 635 152
rect 637 150 640 152
rect 663 152 677 154
rect 663 151 670 152
rect 631 142 640 150
rect 647 142 652 151
rect 631 129 642 142
rect 644 133 652 142
rect 644 131 647 133
rect 649 131 652 133
rect 644 129 652 131
rect 611 127 618 129
rect 647 126 652 129
rect 654 126 659 151
rect 661 150 670 151
rect 672 150 677 152
rect 661 145 677 150
rect 661 143 670 145
rect 672 143 677 145
rect 661 126 677 143
rect 679 144 687 154
rect 679 142 682 144
rect 684 142 687 144
rect 679 137 687 142
rect 679 135 682 137
rect 684 135 687 137
rect 679 126 687 135
rect 689 152 697 154
rect 689 150 692 152
rect 694 150 697 152
rect 689 145 697 150
rect 689 143 692 145
rect 694 143 697 145
rect 689 126 697 143
rect 699 139 704 154
rect 714 139 719 154
rect 699 137 706 139
rect 699 135 702 137
rect 704 135 706 137
rect 699 130 706 135
rect 699 128 702 130
rect 704 128 706 130
rect 699 126 706 128
rect 712 137 719 139
rect 712 135 714 137
rect 716 135 719 137
rect 712 130 719 135
rect 712 128 714 130
rect 716 128 719 130
rect 712 126 719 128
rect 721 152 729 154
rect 721 150 724 152
rect 726 150 729 152
rect 721 145 729 150
rect 721 143 724 145
rect 726 143 729 145
rect 721 126 729 143
rect 731 144 739 154
rect 731 142 734 144
rect 736 142 739 144
rect 731 137 739 142
rect 731 135 734 137
rect 736 135 739 137
rect 731 126 739 135
rect 741 152 755 154
rect 741 150 746 152
rect 748 151 755 152
rect 778 152 787 154
rect 748 150 757 151
rect 741 145 757 150
rect 741 143 746 145
rect 748 143 757 145
rect 741 126 757 143
rect 759 126 764 151
rect 766 142 771 151
rect 778 150 781 152
rect 783 150 787 152
rect 778 142 787 150
rect 766 133 774 142
rect 766 131 769 133
rect 771 131 774 133
rect 766 129 774 131
rect 776 129 787 142
rect 789 142 794 154
rect 803 147 808 154
rect 801 145 808 147
rect 801 143 803 145
rect 805 143 808 145
rect 789 140 796 142
rect 801 141 808 143
rect 789 138 792 140
rect 794 138 796 140
rect 789 133 796 138
rect 803 133 808 141
rect 810 133 815 154
rect 817 152 826 154
rect 817 150 822 152
rect 824 150 826 152
rect 817 144 826 150
rect 849 145 856 147
rect 817 133 828 144
rect 789 131 792 133
rect 794 131 796 133
rect 789 129 796 131
rect 766 126 771 129
rect 820 126 828 133
rect 830 142 837 144
rect 830 140 833 142
rect 835 140 837 142
rect 830 135 837 140
rect 830 133 833 135
rect 835 133 837 135
rect 849 143 851 145
rect 853 143 856 145
rect 849 134 856 143
rect 858 145 866 147
rect 858 143 861 145
rect 863 143 866 145
rect 858 138 866 143
rect 858 136 861 138
rect 863 136 866 138
rect 858 134 866 136
rect 868 145 874 147
rect 868 143 876 145
rect 868 141 871 143
rect 873 141 876 143
rect 868 134 876 141
rect 830 131 837 133
rect 830 126 835 131
rect 870 127 876 134
rect 878 140 883 145
rect 891 142 896 154
rect 889 140 896 142
rect 878 138 885 140
rect 878 136 881 138
rect 883 136 885 138
rect 878 131 885 136
rect 878 129 881 131
rect 883 129 885 131
rect 889 138 891 140
rect 893 138 896 140
rect 889 133 896 138
rect 889 131 891 133
rect 893 131 896 133
rect 889 129 896 131
rect 898 152 907 154
rect 898 150 902 152
rect 904 150 907 152
rect 930 152 944 154
rect 930 151 937 152
rect 898 142 907 150
rect 914 142 919 151
rect 898 129 909 142
rect 911 133 919 142
rect 911 131 914 133
rect 916 131 919 133
rect 911 129 919 131
rect 878 127 885 129
rect 914 126 919 129
rect 921 126 926 151
rect 928 150 937 151
rect 939 150 944 152
rect 928 145 944 150
rect 928 143 937 145
rect 939 143 944 145
rect 928 126 944 143
rect 946 144 954 154
rect 946 142 949 144
rect 951 142 954 144
rect 946 137 954 142
rect 946 135 949 137
rect 951 135 954 137
rect 946 126 954 135
rect 956 152 964 154
rect 956 150 959 152
rect 961 150 964 152
rect 956 145 964 150
rect 956 143 959 145
rect 961 143 964 145
rect 956 126 964 143
rect 966 139 971 154
rect 981 139 986 154
rect 966 137 973 139
rect 966 135 969 137
rect 971 135 973 137
rect 966 130 973 135
rect 966 128 969 130
rect 971 128 973 130
rect 966 126 973 128
rect 979 137 986 139
rect 979 135 981 137
rect 983 135 986 137
rect 979 130 986 135
rect 979 128 981 130
rect 983 128 986 130
rect 979 126 986 128
rect 988 152 996 154
rect 988 150 991 152
rect 993 150 996 152
rect 988 145 996 150
rect 988 143 991 145
rect 993 143 996 145
rect 988 126 996 143
rect 998 144 1006 154
rect 998 142 1001 144
rect 1003 142 1006 144
rect 998 137 1006 142
rect 998 135 1001 137
rect 1003 135 1006 137
rect 998 126 1006 135
rect 1008 152 1022 154
rect 1008 150 1013 152
rect 1015 151 1022 152
rect 1045 152 1054 154
rect 1015 150 1024 151
rect 1008 145 1024 150
rect 1008 143 1013 145
rect 1015 143 1024 145
rect 1008 126 1024 143
rect 1026 126 1031 151
rect 1033 142 1038 151
rect 1045 150 1048 152
rect 1050 150 1054 152
rect 1045 142 1054 150
rect 1033 133 1041 142
rect 1033 131 1036 133
rect 1038 131 1041 133
rect 1033 129 1041 131
rect 1043 129 1054 142
rect 1056 142 1061 154
rect 1070 147 1075 154
rect 1068 145 1075 147
rect 1068 143 1070 145
rect 1072 143 1075 145
rect 1056 140 1063 142
rect 1068 141 1075 143
rect 1056 138 1059 140
rect 1061 138 1063 140
rect 1056 133 1063 138
rect 1070 133 1075 141
rect 1077 133 1082 154
rect 1084 152 1093 154
rect 1084 150 1089 152
rect 1091 150 1093 152
rect 1084 144 1093 150
rect 1116 145 1123 147
rect 1084 133 1095 144
rect 1056 131 1059 133
rect 1061 131 1063 133
rect 1056 129 1063 131
rect 1033 126 1038 129
rect 1087 126 1095 133
rect 1097 142 1104 144
rect 1097 140 1100 142
rect 1102 140 1104 142
rect 1097 135 1104 140
rect 1097 133 1100 135
rect 1102 133 1104 135
rect 1116 143 1118 145
rect 1120 143 1123 145
rect 1116 134 1123 143
rect 1125 145 1133 147
rect 1125 143 1128 145
rect 1130 143 1133 145
rect 1125 138 1133 143
rect 1125 136 1128 138
rect 1130 136 1133 138
rect 1125 134 1133 136
rect 1135 145 1141 147
rect 1135 143 1143 145
rect 1135 141 1138 143
rect 1140 141 1143 143
rect 1135 134 1143 141
rect 1097 131 1104 133
rect 1097 126 1102 131
rect 1137 127 1143 134
rect 1145 140 1150 145
rect 1158 142 1163 154
rect 1156 140 1163 142
rect 1145 138 1152 140
rect 1145 136 1148 138
rect 1150 136 1152 138
rect 1145 131 1152 136
rect 1145 129 1148 131
rect 1150 129 1152 131
rect 1156 138 1158 140
rect 1160 138 1163 140
rect 1156 133 1163 138
rect 1156 131 1158 133
rect 1160 131 1163 133
rect 1156 129 1163 131
rect 1165 152 1174 154
rect 1165 150 1169 152
rect 1171 150 1174 152
rect 1197 152 1211 154
rect 1197 151 1204 152
rect 1165 142 1174 150
rect 1181 142 1186 151
rect 1165 129 1176 142
rect 1178 133 1186 142
rect 1178 131 1181 133
rect 1183 131 1186 133
rect 1178 129 1186 131
rect 1145 127 1152 129
rect 1181 126 1186 129
rect 1188 126 1193 151
rect 1195 150 1204 151
rect 1206 150 1211 152
rect 1195 145 1211 150
rect 1195 143 1204 145
rect 1206 143 1211 145
rect 1195 126 1211 143
rect 1213 144 1221 154
rect 1213 142 1216 144
rect 1218 142 1221 144
rect 1213 137 1221 142
rect 1213 135 1216 137
rect 1218 135 1221 137
rect 1213 126 1221 135
rect 1223 152 1231 154
rect 1223 150 1226 152
rect 1228 150 1231 152
rect 1223 145 1231 150
rect 1223 143 1226 145
rect 1228 143 1231 145
rect 1223 126 1231 143
rect 1233 139 1238 154
rect 1248 139 1253 154
rect 1233 137 1240 139
rect 1233 135 1236 137
rect 1238 135 1240 137
rect 1233 130 1240 135
rect 1233 128 1236 130
rect 1238 128 1240 130
rect 1233 126 1240 128
rect 1246 137 1253 139
rect 1246 135 1248 137
rect 1250 135 1253 137
rect 1246 130 1253 135
rect 1246 128 1248 130
rect 1250 128 1253 130
rect 1246 126 1253 128
rect 1255 152 1263 154
rect 1255 150 1258 152
rect 1260 150 1263 152
rect 1255 145 1263 150
rect 1255 143 1258 145
rect 1260 143 1263 145
rect 1255 126 1263 143
rect 1265 144 1273 154
rect 1265 142 1268 144
rect 1270 142 1273 144
rect 1265 137 1273 142
rect 1265 135 1268 137
rect 1270 135 1273 137
rect 1265 126 1273 135
rect 1275 152 1289 154
rect 1275 150 1280 152
rect 1282 151 1289 152
rect 1312 152 1321 154
rect 1282 150 1291 151
rect 1275 145 1291 150
rect 1275 143 1280 145
rect 1282 143 1291 145
rect 1275 126 1291 143
rect 1293 126 1298 151
rect 1300 142 1305 151
rect 1312 150 1315 152
rect 1317 150 1321 152
rect 1312 142 1321 150
rect 1300 133 1308 142
rect 1300 131 1303 133
rect 1305 131 1308 133
rect 1300 129 1308 131
rect 1310 129 1321 142
rect 1323 142 1328 154
rect 1337 147 1342 154
rect 1335 145 1342 147
rect 1335 143 1337 145
rect 1339 143 1342 145
rect 1323 140 1330 142
rect 1335 141 1342 143
rect 1323 138 1326 140
rect 1328 138 1330 140
rect 1323 133 1330 138
rect 1337 133 1342 141
rect 1344 133 1349 154
rect 1351 152 1360 154
rect 1351 150 1356 152
rect 1358 150 1360 152
rect 1351 144 1360 150
rect 1383 145 1390 147
rect 1351 133 1362 144
rect 1323 131 1326 133
rect 1328 131 1330 133
rect 1323 129 1330 131
rect 1300 126 1305 129
rect 1354 126 1362 133
rect 1364 142 1371 144
rect 1364 140 1367 142
rect 1369 140 1371 142
rect 1364 135 1371 140
rect 1364 133 1367 135
rect 1369 133 1371 135
rect 1383 143 1385 145
rect 1387 143 1390 145
rect 1383 134 1390 143
rect 1392 145 1400 147
rect 1392 143 1395 145
rect 1397 143 1400 145
rect 1392 138 1400 143
rect 1392 136 1395 138
rect 1397 136 1400 138
rect 1392 134 1400 136
rect 1402 145 1408 147
rect 1402 143 1410 145
rect 1402 141 1405 143
rect 1407 141 1410 143
rect 1402 134 1410 141
rect 1364 131 1371 133
rect 1364 126 1369 131
rect 1404 127 1410 134
rect 1412 140 1417 145
rect 1425 142 1430 154
rect 1423 140 1430 142
rect 1412 138 1419 140
rect 1412 136 1415 138
rect 1417 136 1419 138
rect 1412 131 1419 136
rect 1412 129 1415 131
rect 1417 129 1419 131
rect 1423 138 1425 140
rect 1427 138 1430 140
rect 1423 133 1430 138
rect 1423 131 1425 133
rect 1427 131 1430 133
rect 1423 129 1430 131
rect 1432 152 1441 154
rect 1432 150 1436 152
rect 1438 150 1441 152
rect 1464 152 1478 154
rect 1464 151 1471 152
rect 1432 142 1441 150
rect 1448 142 1453 151
rect 1432 129 1443 142
rect 1445 133 1453 142
rect 1445 131 1448 133
rect 1450 131 1453 133
rect 1445 129 1453 131
rect 1412 127 1419 129
rect 1448 126 1453 129
rect 1455 126 1460 151
rect 1462 150 1471 151
rect 1473 150 1478 152
rect 1462 145 1478 150
rect 1462 143 1471 145
rect 1473 143 1478 145
rect 1462 126 1478 143
rect 1480 144 1488 154
rect 1480 142 1483 144
rect 1485 142 1488 144
rect 1480 137 1488 142
rect 1480 135 1483 137
rect 1485 135 1488 137
rect 1480 126 1488 135
rect 1490 152 1498 154
rect 1490 150 1493 152
rect 1495 150 1498 152
rect 1490 145 1498 150
rect 1490 143 1493 145
rect 1495 143 1498 145
rect 1490 126 1498 143
rect 1500 139 1505 154
rect 1515 139 1520 154
rect 1500 137 1507 139
rect 1500 135 1503 137
rect 1505 135 1507 137
rect 1500 130 1507 135
rect 1500 128 1503 130
rect 1505 128 1507 130
rect 1500 126 1507 128
rect 1513 137 1520 139
rect 1513 135 1515 137
rect 1517 135 1520 137
rect 1513 130 1520 135
rect 1513 128 1515 130
rect 1517 128 1520 130
rect 1513 126 1520 128
rect 1522 152 1530 154
rect 1522 150 1525 152
rect 1527 150 1530 152
rect 1522 145 1530 150
rect 1522 143 1525 145
rect 1527 143 1530 145
rect 1522 126 1530 143
rect 1532 144 1540 154
rect 1532 142 1535 144
rect 1537 142 1540 144
rect 1532 137 1540 142
rect 1532 135 1535 137
rect 1537 135 1540 137
rect 1532 126 1540 135
rect 1542 152 1556 154
rect 1542 150 1547 152
rect 1549 151 1556 152
rect 1579 152 1588 154
rect 1549 150 1558 151
rect 1542 145 1558 150
rect 1542 143 1547 145
rect 1549 143 1558 145
rect 1542 126 1558 143
rect 1560 126 1565 151
rect 1567 142 1572 151
rect 1579 150 1582 152
rect 1584 150 1588 152
rect 1579 142 1588 150
rect 1567 133 1575 142
rect 1567 131 1570 133
rect 1572 131 1575 133
rect 1567 129 1575 131
rect 1577 129 1588 142
rect 1590 142 1595 154
rect 1604 147 1609 154
rect 1602 145 1609 147
rect 1602 143 1604 145
rect 1606 143 1609 145
rect 1590 140 1597 142
rect 1602 141 1609 143
rect 1590 138 1593 140
rect 1595 138 1597 140
rect 1590 133 1597 138
rect 1604 133 1609 141
rect 1611 133 1616 154
rect 1618 152 1627 154
rect 1618 150 1623 152
rect 1625 150 1627 152
rect 1618 144 1627 150
rect 1650 145 1657 147
rect 1618 133 1629 144
rect 1590 131 1593 133
rect 1595 131 1597 133
rect 1590 129 1597 131
rect 1567 126 1572 129
rect 1621 126 1629 133
rect 1631 142 1638 144
rect 1631 140 1634 142
rect 1636 140 1638 142
rect 1631 135 1638 140
rect 1631 133 1634 135
rect 1636 133 1638 135
rect 1650 143 1652 145
rect 1654 143 1657 145
rect 1650 134 1657 143
rect 1659 145 1667 147
rect 1659 143 1662 145
rect 1664 143 1667 145
rect 1659 138 1667 143
rect 1659 136 1662 138
rect 1664 136 1667 138
rect 1659 134 1667 136
rect 1669 145 1675 147
rect 1669 143 1677 145
rect 1669 141 1672 143
rect 1674 141 1677 143
rect 1669 134 1677 141
rect 1631 131 1638 133
rect 1631 126 1636 131
rect 1671 127 1677 134
rect 1679 140 1684 145
rect 1692 142 1697 154
rect 1690 140 1697 142
rect 1679 138 1686 140
rect 1679 136 1682 138
rect 1684 136 1686 138
rect 1679 131 1686 136
rect 1679 129 1682 131
rect 1684 129 1686 131
rect 1690 138 1692 140
rect 1694 138 1697 140
rect 1690 133 1697 138
rect 1690 131 1692 133
rect 1694 131 1697 133
rect 1690 129 1697 131
rect 1699 152 1708 154
rect 1699 150 1703 152
rect 1705 150 1708 152
rect 1731 152 1745 154
rect 1731 151 1738 152
rect 1699 142 1708 150
rect 1715 142 1720 151
rect 1699 129 1710 142
rect 1712 133 1720 142
rect 1712 131 1715 133
rect 1717 131 1720 133
rect 1712 129 1720 131
rect 1679 127 1686 129
rect 1715 126 1720 129
rect 1722 126 1727 151
rect 1729 150 1738 151
rect 1740 150 1745 152
rect 1729 145 1745 150
rect 1729 143 1738 145
rect 1740 143 1745 145
rect 1729 126 1745 143
rect 1747 144 1755 154
rect 1747 142 1750 144
rect 1752 142 1755 144
rect 1747 137 1755 142
rect 1747 135 1750 137
rect 1752 135 1755 137
rect 1747 126 1755 135
rect 1757 152 1765 154
rect 1757 150 1760 152
rect 1762 150 1765 152
rect 1757 145 1765 150
rect 1757 143 1760 145
rect 1762 143 1765 145
rect 1757 126 1765 143
rect 1767 139 1772 154
rect 1782 139 1787 154
rect 1767 137 1774 139
rect 1767 135 1770 137
rect 1772 135 1774 137
rect 1767 130 1774 135
rect 1767 128 1770 130
rect 1772 128 1774 130
rect 1767 126 1774 128
rect 1780 137 1787 139
rect 1780 135 1782 137
rect 1784 135 1787 137
rect 1780 130 1787 135
rect 1780 128 1782 130
rect 1784 128 1787 130
rect 1780 126 1787 128
rect 1789 152 1797 154
rect 1789 150 1792 152
rect 1794 150 1797 152
rect 1789 145 1797 150
rect 1789 143 1792 145
rect 1794 143 1797 145
rect 1789 126 1797 143
rect 1799 144 1807 154
rect 1799 142 1802 144
rect 1804 142 1807 144
rect 1799 137 1807 142
rect 1799 135 1802 137
rect 1804 135 1807 137
rect 1799 126 1807 135
rect 1809 152 1823 154
rect 1809 150 1814 152
rect 1816 151 1823 152
rect 1846 152 1855 154
rect 1816 150 1825 151
rect 1809 145 1825 150
rect 1809 143 1814 145
rect 1816 143 1825 145
rect 1809 126 1825 143
rect 1827 126 1832 151
rect 1834 142 1839 151
rect 1846 150 1849 152
rect 1851 150 1855 152
rect 1846 142 1855 150
rect 1834 133 1842 142
rect 1834 131 1837 133
rect 1839 131 1842 133
rect 1834 129 1842 131
rect 1844 129 1855 142
rect 1857 142 1862 154
rect 1871 147 1876 154
rect 1869 145 1876 147
rect 1869 143 1871 145
rect 1873 143 1876 145
rect 1857 140 1864 142
rect 1869 141 1876 143
rect 1857 138 1860 140
rect 1862 138 1864 140
rect 1857 133 1864 138
rect 1871 133 1876 141
rect 1878 133 1883 154
rect 1885 152 1894 154
rect 1885 150 1890 152
rect 1892 150 1894 152
rect 1885 144 1894 150
rect 1885 133 1896 144
rect 1857 131 1860 133
rect 1862 131 1864 133
rect 1857 129 1864 131
rect 1834 126 1839 129
rect 1888 126 1896 133
rect 1898 142 1905 144
rect 1898 140 1901 142
rect 1903 140 1905 142
rect 1898 135 1905 140
rect 1898 133 1901 135
rect 1903 133 1905 135
rect 1922 133 1927 154
rect 1898 131 1905 133
rect 1920 131 1927 133
rect 1898 126 1903 131
rect 1920 129 1922 131
rect 1924 129 1927 131
rect 1920 127 1927 129
rect 1929 152 1941 154
rect 1929 150 1932 152
rect 1934 150 1941 152
rect 1929 145 1941 150
rect 1958 145 1963 154
rect 1929 143 1932 145
rect 1934 143 1943 145
rect 1929 127 1943 143
rect 1945 138 1953 145
rect 1945 136 1948 138
rect 1950 136 1953 138
rect 1945 131 1953 136
rect 1945 129 1948 131
rect 1950 129 1953 131
rect 1945 127 1953 129
rect 1955 138 1963 145
rect 1955 136 1958 138
rect 1960 136 1963 138
rect 1955 127 1963 136
rect 1965 148 1970 154
rect 1965 146 1972 148
rect 1965 144 1968 146
rect 1970 144 1972 146
rect 1965 142 1972 144
rect 1978 142 1983 154
rect 1965 127 1970 142
rect 1976 140 1983 142
rect 1976 138 1978 140
rect 1980 138 1983 140
rect 1976 133 1983 138
rect 1976 131 1978 133
rect 1980 131 1983 133
rect 1976 129 1983 131
rect 1985 152 1994 154
rect 1985 150 1989 152
rect 1991 150 1994 152
rect 2017 152 2031 154
rect 2017 151 2024 152
rect 1985 142 1994 150
rect 2001 142 2006 151
rect 1985 129 1996 142
rect 1998 133 2006 142
rect 1998 131 2001 133
rect 2003 131 2006 133
rect 1998 129 2006 131
rect 2001 126 2006 129
rect 2008 126 2013 151
rect 2015 150 2024 151
rect 2026 150 2031 152
rect 2015 145 2031 150
rect 2015 143 2024 145
rect 2026 143 2031 145
rect 2015 126 2031 143
rect 2033 144 2041 154
rect 2033 142 2036 144
rect 2038 142 2041 144
rect 2033 137 2041 142
rect 2033 135 2036 137
rect 2038 135 2041 137
rect 2033 126 2041 135
rect 2043 152 2051 154
rect 2043 150 2046 152
rect 2048 150 2051 152
rect 2043 145 2051 150
rect 2043 143 2046 145
rect 2048 143 2051 145
rect 2043 126 2051 143
rect 2053 139 2058 154
rect 2068 139 2073 154
rect 2053 137 2060 139
rect 2053 135 2056 137
rect 2058 135 2060 137
rect 2053 130 2060 135
rect 2053 128 2056 130
rect 2058 128 2060 130
rect 2053 126 2060 128
rect 2066 137 2073 139
rect 2066 135 2068 137
rect 2070 135 2073 137
rect 2066 130 2073 135
rect 2066 128 2068 130
rect 2070 128 2073 130
rect 2066 126 2073 128
rect 2075 152 2083 154
rect 2075 150 2078 152
rect 2080 150 2083 152
rect 2075 145 2083 150
rect 2075 143 2078 145
rect 2080 143 2083 145
rect 2075 126 2083 143
rect 2085 144 2093 154
rect 2085 142 2088 144
rect 2090 142 2093 144
rect 2085 137 2093 142
rect 2085 135 2088 137
rect 2090 135 2093 137
rect 2085 126 2093 135
rect 2095 152 2109 154
rect 2095 150 2100 152
rect 2102 151 2109 152
rect 2132 152 2141 154
rect 2102 150 2111 151
rect 2095 145 2111 150
rect 2095 143 2100 145
rect 2102 143 2111 145
rect 2095 126 2111 143
rect 2113 126 2118 151
rect 2120 142 2125 151
rect 2132 150 2135 152
rect 2137 150 2141 152
rect 2132 142 2141 150
rect 2120 133 2128 142
rect 2120 131 2123 133
rect 2125 131 2128 133
rect 2120 129 2128 131
rect 2130 129 2141 142
rect 2143 142 2148 154
rect 2157 147 2162 154
rect 2155 145 2162 147
rect 2155 143 2157 145
rect 2159 143 2162 145
rect 2143 140 2150 142
rect 2155 141 2162 143
rect 2143 138 2146 140
rect 2148 138 2150 140
rect 2143 133 2150 138
rect 2157 133 2162 141
rect 2164 133 2169 154
rect 2171 152 2180 154
rect 2171 150 2176 152
rect 2178 150 2180 152
rect 2209 152 2216 154
rect 2171 144 2180 150
rect 2209 150 2211 152
rect 2213 150 2216 152
rect 2171 133 2182 144
rect 2143 131 2146 133
rect 2148 131 2150 133
rect 2143 129 2150 131
rect 2120 126 2125 129
rect 2174 126 2182 133
rect 2184 142 2191 144
rect 2184 140 2187 142
rect 2189 140 2191 142
rect 2184 135 2191 140
rect 2209 142 2216 150
rect 2184 133 2187 135
rect 2189 133 2191 135
rect 2210 138 2216 142
rect 2218 138 2223 154
rect 2225 142 2233 154
rect 2225 140 2228 142
rect 2230 140 2233 142
rect 2225 138 2233 140
rect 2235 138 2240 154
rect 2242 152 2250 154
rect 2242 150 2245 152
rect 2247 150 2250 152
rect 2242 138 2250 150
rect 2210 134 2214 138
rect 2184 131 2191 133
rect 2201 132 2206 134
rect 2184 126 2189 131
rect 2199 130 2206 132
rect 2199 128 2201 130
rect 2203 128 2206 130
rect 2199 126 2206 128
rect 2208 126 2214 134
rect 2245 136 2250 138
rect 2252 147 2257 154
rect 2277 152 2284 154
rect 2277 150 2279 152
rect 2281 150 2284 152
rect 2252 145 2259 147
rect 2252 143 2255 145
rect 2257 143 2259 145
rect 2252 141 2259 143
rect 2277 142 2284 150
rect 2252 136 2257 141
rect 2278 138 2284 142
rect 2286 138 2291 154
rect 2293 142 2301 154
rect 2293 140 2296 142
rect 2298 140 2301 142
rect 2293 138 2301 140
rect 2303 138 2308 154
rect 2310 152 2318 154
rect 2310 150 2313 152
rect 2315 150 2318 152
rect 2310 138 2318 150
rect 2278 134 2282 138
rect 2269 132 2274 134
rect 2267 130 2274 132
rect 2267 128 2269 130
rect 2271 128 2274 130
rect 2267 126 2274 128
rect 2276 126 2282 134
rect 2313 136 2318 138
rect 2320 147 2325 154
rect 2320 145 2327 147
rect 2320 143 2323 145
rect 2325 143 2327 145
rect 2320 141 2327 143
rect 2320 136 2325 141
rect 29 42 35 49
rect 8 33 15 42
rect 8 31 10 33
rect 12 31 15 33
rect 8 29 15 31
rect 17 40 25 42
rect 17 38 20 40
rect 22 38 25 40
rect 17 33 25 38
rect 17 31 20 33
rect 22 31 25 33
rect 17 29 25 31
rect 27 35 35 42
rect 27 33 30 35
rect 32 33 35 35
rect 27 31 35 33
rect 37 44 44 49
rect 37 42 40 44
rect 42 42 44 44
rect 69 42 75 49
rect 37 37 44 42
rect 37 35 40 37
rect 42 35 44 37
rect 37 33 44 35
rect 48 33 55 42
rect 37 31 42 33
rect 48 31 50 33
rect 52 31 55 33
rect 27 29 33 31
rect 48 29 55 31
rect 57 40 65 42
rect 57 38 60 40
rect 62 38 65 40
rect 57 33 65 38
rect 57 31 60 33
rect 62 31 65 33
rect 57 29 65 31
rect 67 35 75 42
rect 67 33 70 35
rect 72 33 75 35
rect 67 31 75 33
rect 77 47 84 49
rect 113 47 118 50
rect 77 45 80 47
rect 82 45 84 47
rect 77 40 84 45
rect 77 38 80 40
rect 82 38 84 40
rect 77 36 84 38
rect 88 45 95 47
rect 88 43 90 45
rect 92 43 95 45
rect 88 38 95 43
rect 88 36 90 38
rect 92 36 95 38
rect 77 31 82 36
rect 88 34 95 36
rect 67 29 73 31
rect 90 22 95 34
rect 97 34 108 47
rect 110 45 118 47
rect 110 43 113 45
rect 115 43 118 45
rect 110 34 118 43
rect 97 26 106 34
rect 97 24 101 26
rect 103 24 106 26
rect 113 25 118 34
rect 120 25 125 50
rect 127 33 143 50
rect 127 31 136 33
rect 138 31 143 33
rect 127 26 143 31
rect 127 25 136 26
rect 97 22 106 24
rect 129 24 136 25
rect 138 24 143 26
rect 129 22 143 24
rect 145 41 153 50
rect 145 39 148 41
rect 150 39 153 41
rect 145 34 153 39
rect 145 32 148 34
rect 150 32 153 34
rect 145 22 153 32
rect 155 33 163 50
rect 155 31 158 33
rect 160 31 163 33
rect 155 26 163 31
rect 155 24 158 26
rect 160 24 163 26
rect 155 22 163 24
rect 165 48 172 50
rect 165 46 168 48
rect 170 46 172 48
rect 165 41 172 46
rect 165 39 168 41
rect 170 39 172 41
rect 165 37 172 39
rect 178 48 185 50
rect 178 46 180 48
rect 182 46 185 48
rect 178 41 185 46
rect 178 39 180 41
rect 182 39 185 41
rect 178 37 185 39
rect 165 22 170 37
rect 180 22 185 37
rect 187 33 195 50
rect 187 31 190 33
rect 192 31 195 33
rect 187 26 195 31
rect 187 24 190 26
rect 192 24 195 26
rect 187 22 195 24
rect 197 41 205 50
rect 197 39 200 41
rect 202 39 205 41
rect 197 34 205 39
rect 197 32 200 34
rect 202 32 205 34
rect 197 22 205 32
rect 207 33 223 50
rect 207 31 212 33
rect 214 31 223 33
rect 207 26 223 31
rect 207 24 212 26
rect 214 25 223 26
rect 225 25 230 50
rect 232 47 237 50
rect 232 45 240 47
rect 232 43 235 45
rect 237 43 240 45
rect 232 34 240 43
rect 242 34 253 47
rect 232 25 237 34
rect 244 26 253 34
rect 214 24 221 25
rect 207 22 221 24
rect 244 24 247 26
rect 249 24 253 26
rect 244 22 253 24
rect 255 45 262 47
rect 255 43 258 45
rect 260 43 262 45
rect 286 43 294 50
rect 255 38 262 43
rect 255 36 258 38
rect 260 36 262 38
rect 255 34 262 36
rect 269 35 274 43
rect 255 22 260 34
rect 267 33 274 35
rect 267 31 269 33
rect 271 31 274 33
rect 267 29 274 31
rect 269 22 274 29
rect 276 22 281 43
rect 283 32 294 43
rect 296 45 301 50
rect 296 43 303 45
rect 296 41 299 43
rect 301 41 303 43
rect 336 42 342 49
rect 296 36 303 41
rect 296 34 299 36
rect 301 34 303 36
rect 296 32 303 34
rect 315 33 322 42
rect 283 26 292 32
rect 315 31 317 33
rect 319 31 322 33
rect 315 29 322 31
rect 324 40 332 42
rect 324 38 327 40
rect 329 38 332 40
rect 324 33 332 38
rect 324 31 327 33
rect 329 31 332 33
rect 324 29 332 31
rect 334 35 342 42
rect 334 33 337 35
rect 339 33 342 35
rect 334 31 342 33
rect 344 47 351 49
rect 380 47 385 50
rect 344 45 347 47
rect 349 45 351 47
rect 344 40 351 45
rect 344 38 347 40
rect 349 38 351 40
rect 344 36 351 38
rect 355 45 362 47
rect 355 43 357 45
rect 359 43 362 45
rect 355 38 362 43
rect 355 36 357 38
rect 359 36 362 38
rect 344 31 349 36
rect 355 34 362 36
rect 334 29 340 31
rect 283 24 288 26
rect 290 24 292 26
rect 283 22 292 24
rect 357 22 362 34
rect 364 34 375 47
rect 377 45 385 47
rect 377 43 380 45
rect 382 43 385 45
rect 377 34 385 43
rect 364 26 373 34
rect 364 24 368 26
rect 370 24 373 26
rect 380 25 385 34
rect 387 25 392 50
rect 394 33 410 50
rect 394 31 403 33
rect 405 31 410 33
rect 394 26 410 31
rect 394 25 403 26
rect 364 22 373 24
rect 396 24 403 25
rect 405 24 410 26
rect 396 22 410 24
rect 412 41 420 50
rect 412 39 415 41
rect 417 39 420 41
rect 412 34 420 39
rect 412 32 415 34
rect 417 32 420 34
rect 412 22 420 32
rect 422 33 430 50
rect 422 31 425 33
rect 427 31 430 33
rect 422 26 430 31
rect 422 24 425 26
rect 427 24 430 26
rect 422 22 430 24
rect 432 48 439 50
rect 432 46 435 48
rect 437 46 439 48
rect 432 41 439 46
rect 432 39 435 41
rect 437 39 439 41
rect 432 37 439 39
rect 445 48 452 50
rect 445 46 447 48
rect 449 46 452 48
rect 445 41 452 46
rect 445 39 447 41
rect 449 39 452 41
rect 445 37 452 39
rect 432 22 437 37
rect 447 22 452 37
rect 454 33 462 50
rect 454 31 457 33
rect 459 31 462 33
rect 454 26 462 31
rect 454 24 457 26
rect 459 24 462 26
rect 454 22 462 24
rect 464 41 472 50
rect 464 39 467 41
rect 469 39 472 41
rect 464 34 472 39
rect 464 32 467 34
rect 469 32 472 34
rect 464 22 472 32
rect 474 33 490 50
rect 474 31 479 33
rect 481 31 490 33
rect 474 26 490 31
rect 474 24 479 26
rect 481 25 490 26
rect 492 25 497 50
rect 499 47 504 50
rect 499 45 507 47
rect 499 43 502 45
rect 504 43 507 45
rect 499 34 507 43
rect 509 34 520 47
rect 499 25 504 34
rect 511 26 520 34
rect 481 24 488 25
rect 474 22 488 24
rect 511 24 514 26
rect 516 24 520 26
rect 511 22 520 24
rect 522 45 529 47
rect 522 43 525 45
rect 527 43 529 45
rect 553 43 561 50
rect 522 38 529 43
rect 522 36 525 38
rect 527 36 529 38
rect 522 34 529 36
rect 536 35 541 43
rect 522 22 527 34
rect 534 33 541 35
rect 534 31 536 33
rect 538 31 541 33
rect 534 29 541 31
rect 536 22 541 29
rect 543 22 548 43
rect 550 32 561 43
rect 563 45 568 50
rect 563 43 570 45
rect 563 41 566 43
rect 568 41 570 43
rect 603 42 609 49
rect 563 36 570 41
rect 563 34 566 36
rect 568 34 570 36
rect 563 32 570 34
rect 582 33 589 42
rect 550 26 559 32
rect 582 31 584 33
rect 586 31 589 33
rect 582 29 589 31
rect 591 40 599 42
rect 591 38 594 40
rect 596 38 599 40
rect 591 33 599 38
rect 591 31 594 33
rect 596 31 599 33
rect 591 29 599 31
rect 601 35 609 42
rect 601 33 604 35
rect 606 33 609 35
rect 601 31 609 33
rect 611 47 618 49
rect 647 47 652 50
rect 611 45 614 47
rect 616 45 618 47
rect 611 40 618 45
rect 611 38 614 40
rect 616 38 618 40
rect 611 36 618 38
rect 622 45 629 47
rect 622 43 624 45
rect 626 43 629 45
rect 622 38 629 43
rect 622 36 624 38
rect 626 36 629 38
rect 611 31 616 36
rect 622 34 629 36
rect 601 29 607 31
rect 550 24 555 26
rect 557 24 559 26
rect 550 22 559 24
rect 624 22 629 34
rect 631 34 642 47
rect 644 45 652 47
rect 644 43 647 45
rect 649 43 652 45
rect 644 34 652 43
rect 631 26 640 34
rect 631 24 635 26
rect 637 24 640 26
rect 647 25 652 34
rect 654 25 659 50
rect 661 33 677 50
rect 661 31 670 33
rect 672 31 677 33
rect 661 26 677 31
rect 661 25 670 26
rect 631 22 640 24
rect 663 24 670 25
rect 672 24 677 26
rect 663 22 677 24
rect 679 41 687 50
rect 679 39 682 41
rect 684 39 687 41
rect 679 34 687 39
rect 679 32 682 34
rect 684 32 687 34
rect 679 22 687 32
rect 689 33 697 50
rect 689 31 692 33
rect 694 31 697 33
rect 689 26 697 31
rect 689 24 692 26
rect 694 24 697 26
rect 689 22 697 24
rect 699 48 706 50
rect 699 46 702 48
rect 704 46 706 48
rect 699 41 706 46
rect 699 39 702 41
rect 704 39 706 41
rect 699 37 706 39
rect 712 48 719 50
rect 712 46 714 48
rect 716 46 719 48
rect 712 41 719 46
rect 712 39 714 41
rect 716 39 719 41
rect 712 37 719 39
rect 699 22 704 37
rect 714 22 719 37
rect 721 33 729 50
rect 721 31 724 33
rect 726 31 729 33
rect 721 26 729 31
rect 721 24 724 26
rect 726 24 729 26
rect 721 22 729 24
rect 731 41 739 50
rect 731 39 734 41
rect 736 39 739 41
rect 731 34 739 39
rect 731 32 734 34
rect 736 32 739 34
rect 731 22 739 32
rect 741 33 757 50
rect 741 31 746 33
rect 748 31 757 33
rect 741 26 757 31
rect 741 24 746 26
rect 748 25 757 26
rect 759 25 764 50
rect 766 47 771 50
rect 766 45 774 47
rect 766 43 769 45
rect 771 43 774 45
rect 766 34 774 43
rect 776 34 787 47
rect 766 25 771 34
rect 778 26 787 34
rect 748 24 755 25
rect 741 22 755 24
rect 778 24 781 26
rect 783 24 787 26
rect 778 22 787 24
rect 789 45 796 47
rect 789 43 792 45
rect 794 43 796 45
rect 820 43 828 50
rect 789 38 796 43
rect 789 36 792 38
rect 794 36 796 38
rect 789 34 796 36
rect 803 35 808 43
rect 789 22 794 34
rect 801 33 808 35
rect 801 31 803 33
rect 805 31 808 33
rect 801 29 808 31
rect 803 22 808 29
rect 810 22 815 43
rect 817 32 828 43
rect 830 45 835 50
rect 830 43 837 45
rect 830 41 833 43
rect 835 41 837 43
rect 870 42 876 49
rect 830 36 837 41
rect 830 34 833 36
rect 835 34 837 36
rect 830 32 837 34
rect 849 33 856 42
rect 817 26 826 32
rect 849 31 851 33
rect 853 31 856 33
rect 849 29 856 31
rect 858 40 866 42
rect 858 38 861 40
rect 863 38 866 40
rect 858 33 866 38
rect 858 31 861 33
rect 863 31 866 33
rect 858 29 866 31
rect 868 35 876 42
rect 868 33 871 35
rect 873 33 876 35
rect 868 31 876 33
rect 878 47 885 49
rect 914 47 919 50
rect 878 45 881 47
rect 883 45 885 47
rect 878 40 885 45
rect 878 38 881 40
rect 883 38 885 40
rect 878 36 885 38
rect 889 45 896 47
rect 889 43 891 45
rect 893 43 896 45
rect 889 38 896 43
rect 889 36 891 38
rect 893 36 896 38
rect 878 31 883 36
rect 889 34 896 36
rect 868 29 874 31
rect 817 24 822 26
rect 824 24 826 26
rect 817 22 826 24
rect 891 22 896 34
rect 898 34 909 47
rect 911 45 919 47
rect 911 43 914 45
rect 916 43 919 45
rect 911 34 919 43
rect 898 26 907 34
rect 898 24 902 26
rect 904 24 907 26
rect 914 25 919 34
rect 921 25 926 50
rect 928 33 944 50
rect 928 31 937 33
rect 939 31 944 33
rect 928 26 944 31
rect 928 25 937 26
rect 898 22 907 24
rect 930 24 937 25
rect 939 24 944 26
rect 930 22 944 24
rect 946 41 954 50
rect 946 39 949 41
rect 951 39 954 41
rect 946 34 954 39
rect 946 32 949 34
rect 951 32 954 34
rect 946 22 954 32
rect 956 33 964 50
rect 956 31 959 33
rect 961 31 964 33
rect 956 26 964 31
rect 956 24 959 26
rect 961 24 964 26
rect 956 22 964 24
rect 966 48 973 50
rect 966 46 969 48
rect 971 46 973 48
rect 966 41 973 46
rect 966 39 969 41
rect 971 39 973 41
rect 966 37 973 39
rect 979 48 986 50
rect 979 46 981 48
rect 983 46 986 48
rect 979 41 986 46
rect 979 39 981 41
rect 983 39 986 41
rect 979 37 986 39
rect 966 22 971 37
rect 981 22 986 37
rect 988 33 996 50
rect 988 31 991 33
rect 993 31 996 33
rect 988 26 996 31
rect 988 24 991 26
rect 993 24 996 26
rect 988 22 996 24
rect 998 41 1006 50
rect 998 39 1001 41
rect 1003 39 1006 41
rect 998 34 1006 39
rect 998 32 1001 34
rect 1003 32 1006 34
rect 998 22 1006 32
rect 1008 33 1024 50
rect 1008 31 1013 33
rect 1015 31 1024 33
rect 1008 26 1024 31
rect 1008 24 1013 26
rect 1015 25 1024 26
rect 1026 25 1031 50
rect 1033 47 1038 50
rect 1033 45 1041 47
rect 1033 43 1036 45
rect 1038 43 1041 45
rect 1033 34 1041 43
rect 1043 34 1054 47
rect 1033 25 1038 34
rect 1045 26 1054 34
rect 1015 24 1022 25
rect 1008 22 1022 24
rect 1045 24 1048 26
rect 1050 24 1054 26
rect 1045 22 1054 24
rect 1056 45 1063 47
rect 1056 43 1059 45
rect 1061 43 1063 45
rect 1087 43 1095 50
rect 1056 38 1063 43
rect 1056 36 1059 38
rect 1061 36 1063 38
rect 1056 34 1063 36
rect 1070 35 1075 43
rect 1056 22 1061 34
rect 1068 33 1075 35
rect 1068 31 1070 33
rect 1072 31 1075 33
rect 1068 29 1075 31
rect 1070 22 1075 29
rect 1077 22 1082 43
rect 1084 32 1095 43
rect 1097 45 1102 50
rect 1097 43 1104 45
rect 1097 41 1100 43
rect 1102 41 1104 43
rect 1137 42 1143 49
rect 1097 36 1104 41
rect 1097 34 1100 36
rect 1102 34 1104 36
rect 1097 32 1104 34
rect 1116 33 1123 42
rect 1084 26 1093 32
rect 1116 31 1118 33
rect 1120 31 1123 33
rect 1116 29 1123 31
rect 1125 40 1133 42
rect 1125 38 1128 40
rect 1130 38 1133 40
rect 1125 33 1133 38
rect 1125 31 1128 33
rect 1130 31 1133 33
rect 1125 29 1133 31
rect 1135 35 1143 42
rect 1135 33 1138 35
rect 1140 33 1143 35
rect 1135 31 1143 33
rect 1145 47 1152 49
rect 1181 47 1186 50
rect 1145 45 1148 47
rect 1150 45 1152 47
rect 1145 40 1152 45
rect 1145 38 1148 40
rect 1150 38 1152 40
rect 1145 36 1152 38
rect 1156 45 1163 47
rect 1156 43 1158 45
rect 1160 43 1163 45
rect 1156 38 1163 43
rect 1156 36 1158 38
rect 1160 36 1163 38
rect 1145 31 1150 36
rect 1156 34 1163 36
rect 1135 29 1141 31
rect 1084 24 1089 26
rect 1091 24 1093 26
rect 1084 22 1093 24
rect 1158 22 1163 34
rect 1165 34 1176 47
rect 1178 45 1186 47
rect 1178 43 1181 45
rect 1183 43 1186 45
rect 1178 34 1186 43
rect 1165 26 1174 34
rect 1165 24 1169 26
rect 1171 24 1174 26
rect 1181 25 1186 34
rect 1188 25 1193 50
rect 1195 33 1211 50
rect 1195 31 1204 33
rect 1206 31 1211 33
rect 1195 26 1211 31
rect 1195 25 1204 26
rect 1165 22 1174 24
rect 1197 24 1204 25
rect 1206 24 1211 26
rect 1197 22 1211 24
rect 1213 41 1221 50
rect 1213 39 1216 41
rect 1218 39 1221 41
rect 1213 34 1221 39
rect 1213 32 1216 34
rect 1218 32 1221 34
rect 1213 22 1221 32
rect 1223 33 1231 50
rect 1223 31 1226 33
rect 1228 31 1231 33
rect 1223 26 1231 31
rect 1223 24 1226 26
rect 1228 24 1231 26
rect 1223 22 1231 24
rect 1233 48 1240 50
rect 1233 46 1236 48
rect 1238 46 1240 48
rect 1233 41 1240 46
rect 1233 39 1236 41
rect 1238 39 1240 41
rect 1233 37 1240 39
rect 1246 48 1253 50
rect 1246 46 1248 48
rect 1250 46 1253 48
rect 1246 41 1253 46
rect 1246 39 1248 41
rect 1250 39 1253 41
rect 1246 37 1253 39
rect 1233 22 1238 37
rect 1248 22 1253 37
rect 1255 33 1263 50
rect 1255 31 1258 33
rect 1260 31 1263 33
rect 1255 26 1263 31
rect 1255 24 1258 26
rect 1260 24 1263 26
rect 1255 22 1263 24
rect 1265 41 1273 50
rect 1265 39 1268 41
rect 1270 39 1273 41
rect 1265 34 1273 39
rect 1265 32 1268 34
rect 1270 32 1273 34
rect 1265 22 1273 32
rect 1275 33 1291 50
rect 1275 31 1280 33
rect 1282 31 1291 33
rect 1275 26 1291 31
rect 1275 24 1280 26
rect 1282 25 1291 26
rect 1293 25 1298 50
rect 1300 47 1305 50
rect 1300 45 1308 47
rect 1300 43 1303 45
rect 1305 43 1308 45
rect 1300 34 1308 43
rect 1310 34 1321 47
rect 1300 25 1305 34
rect 1312 26 1321 34
rect 1282 24 1289 25
rect 1275 22 1289 24
rect 1312 24 1315 26
rect 1317 24 1321 26
rect 1312 22 1321 24
rect 1323 45 1330 47
rect 1323 43 1326 45
rect 1328 43 1330 45
rect 1354 43 1362 50
rect 1323 38 1330 43
rect 1323 36 1326 38
rect 1328 36 1330 38
rect 1323 34 1330 36
rect 1337 35 1342 43
rect 1323 22 1328 34
rect 1335 33 1342 35
rect 1335 31 1337 33
rect 1339 31 1342 33
rect 1335 29 1342 31
rect 1337 22 1342 29
rect 1344 22 1349 43
rect 1351 32 1362 43
rect 1364 45 1369 50
rect 1364 43 1371 45
rect 1364 41 1367 43
rect 1369 41 1371 43
rect 1404 42 1410 49
rect 1364 36 1371 41
rect 1364 34 1367 36
rect 1369 34 1371 36
rect 1364 32 1371 34
rect 1383 33 1390 42
rect 1351 26 1360 32
rect 1383 31 1385 33
rect 1387 31 1390 33
rect 1383 29 1390 31
rect 1392 40 1400 42
rect 1392 38 1395 40
rect 1397 38 1400 40
rect 1392 33 1400 38
rect 1392 31 1395 33
rect 1397 31 1400 33
rect 1392 29 1400 31
rect 1402 35 1410 42
rect 1402 33 1405 35
rect 1407 33 1410 35
rect 1402 31 1410 33
rect 1412 47 1419 49
rect 1448 47 1453 50
rect 1412 45 1415 47
rect 1417 45 1419 47
rect 1412 40 1419 45
rect 1412 38 1415 40
rect 1417 38 1419 40
rect 1412 36 1419 38
rect 1423 45 1430 47
rect 1423 43 1425 45
rect 1427 43 1430 45
rect 1423 38 1430 43
rect 1423 36 1425 38
rect 1427 36 1430 38
rect 1412 31 1417 36
rect 1423 34 1430 36
rect 1402 29 1408 31
rect 1351 24 1356 26
rect 1358 24 1360 26
rect 1351 22 1360 24
rect 1425 22 1430 34
rect 1432 34 1443 47
rect 1445 45 1453 47
rect 1445 43 1448 45
rect 1450 43 1453 45
rect 1445 34 1453 43
rect 1432 26 1441 34
rect 1432 24 1436 26
rect 1438 24 1441 26
rect 1448 25 1453 34
rect 1455 25 1460 50
rect 1462 33 1478 50
rect 1462 31 1471 33
rect 1473 31 1478 33
rect 1462 26 1478 31
rect 1462 25 1471 26
rect 1432 22 1441 24
rect 1464 24 1471 25
rect 1473 24 1478 26
rect 1464 22 1478 24
rect 1480 41 1488 50
rect 1480 39 1483 41
rect 1485 39 1488 41
rect 1480 34 1488 39
rect 1480 32 1483 34
rect 1485 32 1488 34
rect 1480 22 1488 32
rect 1490 33 1498 50
rect 1490 31 1493 33
rect 1495 31 1498 33
rect 1490 26 1498 31
rect 1490 24 1493 26
rect 1495 24 1498 26
rect 1490 22 1498 24
rect 1500 48 1507 50
rect 1500 46 1503 48
rect 1505 46 1507 48
rect 1500 41 1507 46
rect 1500 39 1503 41
rect 1505 39 1507 41
rect 1500 37 1507 39
rect 1513 48 1520 50
rect 1513 46 1515 48
rect 1517 46 1520 48
rect 1513 41 1520 46
rect 1513 39 1515 41
rect 1517 39 1520 41
rect 1513 37 1520 39
rect 1500 22 1505 37
rect 1515 22 1520 37
rect 1522 33 1530 50
rect 1522 31 1525 33
rect 1527 31 1530 33
rect 1522 26 1530 31
rect 1522 24 1525 26
rect 1527 24 1530 26
rect 1522 22 1530 24
rect 1532 41 1540 50
rect 1532 39 1535 41
rect 1537 39 1540 41
rect 1532 34 1540 39
rect 1532 32 1535 34
rect 1537 32 1540 34
rect 1532 22 1540 32
rect 1542 33 1558 50
rect 1542 31 1547 33
rect 1549 31 1558 33
rect 1542 26 1558 31
rect 1542 24 1547 26
rect 1549 25 1558 26
rect 1560 25 1565 50
rect 1567 47 1572 50
rect 1567 45 1575 47
rect 1567 43 1570 45
rect 1572 43 1575 45
rect 1567 34 1575 43
rect 1577 34 1588 47
rect 1567 25 1572 34
rect 1579 26 1588 34
rect 1549 24 1556 25
rect 1542 22 1556 24
rect 1579 24 1582 26
rect 1584 24 1588 26
rect 1579 22 1588 24
rect 1590 45 1597 47
rect 1590 43 1593 45
rect 1595 43 1597 45
rect 1621 43 1629 50
rect 1590 38 1597 43
rect 1590 36 1593 38
rect 1595 36 1597 38
rect 1590 34 1597 36
rect 1604 35 1609 43
rect 1590 22 1595 34
rect 1602 33 1609 35
rect 1602 31 1604 33
rect 1606 31 1609 33
rect 1602 29 1609 31
rect 1604 22 1609 29
rect 1611 22 1616 43
rect 1618 32 1629 43
rect 1631 45 1636 50
rect 1631 43 1638 45
rect 1631 41 1634 43
rect 1636 41 1638 43
rect 1671 42 1677 49
rect 1631 36 1638 41
rect 1631 34 1634 36
rect 1636 34 1638 36
rect 1631 32 1638 34
rect 1650 33 1657 42
rect 1618 26 1627 32
rect 1650 31 1652 33
rect 1654 31 1657 33
rect 1650 29 1657 31
rect 1659 40 1667 42
rect 1659 38 1662 40
rect 1664 38 1667 40
rect 1659 33 1667 38
rect 1659 31 1662 33
rect 1664 31 1667 33
rect 1659 29 1667 31
rect 1669 35 1677 42
rect 1669 33 1672 35
rect 1674 33 1677 35
rect 1669 31 1677 33
rect 1679 47 1686 49
rect 1715 47 1720 50
rect 1679 45 1682 47
rect 1684 45 1686 47
rect 1679 40 1686 45
rect 1679 38 1682 40
rect 1684 38 1686 40
rect 1679 36 1686 38
rect 1690 45 1697 47
rect 1690 43 1692 45
rect 1694 43 1697 45
rect 1690 38 1697 43
rect 1690 36 1692 38
rect 1694 36 1697 38
rect 1679 31 1684 36
rect 1690 34 1697 36
rect 1669 29 1675 31
rect 1618 24 1623 26
rect 1625 24 1627 26
rect 1618 22 1627 24
rect 1692 22 1697 34
rect 1699 34 1710 47
rect 1712 45 1720 47
rect 1712 43 1715 45
rect 1717 43 1720 45
rect 1712 34 1720 43
rect 1699 26 1708 34
rect 1699 24 1703 26
rect 1705 24 1708 26
rect 1715 25 1720 34
rect 1722 25 1727 50
rect 1729 33 1745 50
rect 1729 31 1738 33
rect 1740 31 1745 33
rect 1729 26 1745 31
rect 1729 25 1738 26
rect 1699 22 1708 24
rect 1731 24 1738 25
rect 1740 24 1745 26
rect 1731 22 1745 24
rect 1747 41 1755 50
rect 1747 39 1750 41
rect 1752 39 1755 41
rect 1747 34 1755 39
rect 1747 32 1750 34
rect 1752 32 1755 34
rect 1747 22 1755 32
rect 1757 33 1765 50
rect 1757 31 1760 33
rect 1762 31 1765 33
rect 1757 26 1765 31
rect 1757 24 1760 26
rect 1762 24 1765 26
rect 1757 22 1765 24
rect 1767 48 1774 50
rect 1767 46 1770 48
rect 1772 46 1774 48
rect 1767 41 1774 46
rect 1767 39 1770 41
rect 1772 39 1774 41
rect 1767 37 1774 39
rect 1780 48 1787 50
rect 1780 46 1782 48
rect 1784 46 1787 48
rect 1780 41 1787 46
rect 1780 39 1782 41
rect 1784 39 1787 41
rect 1780 37 1787 39
rect 1767 22 1772 37
rect 1782 22 1787 37
rect 1789 33 1797 50
rect 1789 31 1792 33
rect 1794 31 1797 33
rect 1789 26 1797 31
rect 1789 24 1792 26
rect 1794 24 1797 26
rect 1789 22 1797 24
rect 1799 41 1807 50
rect 1799 39 1802 41
rect 1804 39 1807 41
rect 1799 34 1807 39
rect 1799 32 1802 34
rect 1804 32 1807 34
rect 1799 22 1807 32
rect 1809 33 1825 50
rect 1809 31 1814 33
rect 1816 31 1825 33
rect 1809 26 1825 31
rect 1809 24 1814 26
rect 1816 25 1825 26
rect 1827 25 1832 50
rect 1834 47 1839 50
rect 1834 45 1842 47
rect 1834 43 1837 45
rect 1839 43 1842 45
rect 1834 34 1842 43
rect 1844 34 1855 47
rect 1834 25 1839 34
rect 1846 26 1855 34
rect 1816 24 1823 25
rect 1809 22 1823 24
rect 1846 24 1849 26
rect 1851 24 1855 26
rect 1846 22 1855 24
rect 1857 45 1864 47
rect 1857 43 1860 45
rect 1862 43 1864 45
rect 1888 43 1896 50
rect 1857 38 1864 43
rect 1857 36 1860 38
rect 1862 36 1864 38
rect 1857 34 1864 36
rect 1871 35 1876 43
rect 1857 22 1862 34
rect 1869 33 1876 35
rect 1869 31 1871 33
rect 1873 31 1876 33
rect 1869 29 1876 31
rect 1871 22 1876 29
rect 1878 22 1883 43
rect 1885 32 1896 43
rect 1898 45 1903 50
rect 1920 47 1927 49
rect 1920 45 1922 47
rect 1924 45 1927 47
rect 1898 43 1905 45
rect 1920 43 1927 45
rect 1898 41 1901 43
rect 1903 41 1905 43
rect 1898 36 1905 41
rect 1898 34 1901 36
rect 1903 34 1905 36
rect 1898 32 1905 34
rect 1885 26 1894 32
rect 1885 24 1890 26
rect 1892 24 1894 26
rect 1885 22 1894 24
rect 1922 22 1927 43
rect 1929 33 1943 49
rect 1929 31 1932 33
rect 1934 31 1943 33
rect 1945 47 1953 49
rect 1945 45 1948 47
rect 1950 45 1953 47
rect 1945 40 1953 45
rect 1945 38 1948 40
rect 1950 38 1953 40
rect 1945 31 1953 38
rect 1955 40 1963 49
rect 1955 38 1958 40
rect 1960 38 1963 40
rect 1955 31 1963 38
rect 1929 26 1941 31
rect 1929 24 1932 26
rect 1934 24 1941 26
rect 1929 22 1941 24
rect 1958 22 1963 31
rect 1965 34 1970 49
rect 2001 47 2006 50
rect 1976 45 1983 47
rect 1976 43 1978 45
rect 1980 43 1983 45
rect 1976 38 1983 43
rect 1976 36 1978 38
rect 1980 36 1983 38
rect 1976 34 1983 36
rect 1965 32 1972 34
rect 1965 30 1968 32
rect 1970 30 1972 32
rect 1965 28 1972 30
rect 1965 22 1970 28
rect 1978 22 1983 34
rect 1985 34 1996 47
rect 1998 45 2006 47
rect 1998 43 2001 45
rect 2003 43 2006 45
rect 1998 34 2006 43
rect 1985 26 1994 34
rect 1985 24 1989 26
rect 1991 24 1994 26
rect 2001 25 2006 34
rect 2008 25 2013 50
rect 2015 33 2031 50
rect 2015 31 2024 33
rect 2026 31 2031 33
rect 2015 26 2031 31
rect 2015 25 2024 26
rect 1985 22 1994 24
rect 2017 24 2024 25
rect 2026 24 2031 26
rect 2017 22 2031 24
rect 2033 41 2041 50
rect 2033 39 2036 41
rect 2038 39 2041 41
rect 2033 34 2041 39
rect 2033 32 2036 34
rect 2038 32 2041 34
rect 2033 22 2041 32
rect 2043 33 2051 50
rect 2043 31 2046 33
rect 2048 31 2051 33
rect 2043 26 2051 31
rect 2043 24 2046 26
rect 2048 24 2051 26
rect 2043 22 2051 24
rect 2053 48 2060 50
rect 2053 46 2056 48
rect 2058 46 2060 48
rect 2053 41 2060 46
rect 2053 39 2056 41
rect 2058 39 2060 41
rect 2053 37 2060 39
rect 2066 48 2073 50
rect 2066 46 2068 48
rect 2070 46 2073 48
rect 2066 41 2073 46
rect 2066 39 2068 41
rect 2070 39 2073 41
rect 2066 37 2073 39
rect 2053 22 2058 37
rect 2068 22 2073 37
rect 2075 33 2083 50
rect 2075 31 2078 33
rect 2080 31 2083 33
rect 2075 26 2083 31
rect 2075 24 2078 26
rect 2080 24 2083 26
rect 2075 22 2083 24
rect 2085 41 2093 50
rect 2085 39 2088 41
rect 2090 39 2093 41
rect 2085 34 2093 39
rect 2085 32 2088 34
rect 2090 32 2093 34
rect 2085 22 2093 32
rect 2095 33 2111 50
rect 2095 31 2100 33
rect 2102 31 2111 33
rect 2095 26 2111 31
rect 2095 24 2100 26
rect 2102 25 2111 26
rect 2113 25 2118 50
rect 2120 47 2125 50
rect 2120 45 2128 47
rect 2120 43 2123 45
rect 2125 43 2128 45
rect 2120 34 2128 43
rect 2130 34 2141 47
rect 2120 25 2125 34
rect 2132 26 2141 34
rect 2102 24 2109 25
rect 2095 22 2109 24
rect 2132 24 2135 26
rect 2137 24 2141 26
rect 2132 22 2141 24
rect 2143 45 2150 47
rect 2143 43 2146 45
rect 2148 43 2150 45
rect 2174 43 2182 50
rect 2143 38 2150 43
rect 2143 36 2146 38
rect 2148 36 2150 38
rect 2143 34 2150 36
rect 2157 35 2162 43
rect 2143 22 2148 34
rect 2155 33 2162 35
rect 2155 31 2157 33
rect 2159 31 2162 33
rect 2155 29 2162 31
rect 2157 22 2162 29
rect 2164 22 2169 43
rect 2171 32 2182 43
rect 2184 45 2189 50
rect 2199 48 2206 50
rect 2199 46 2201 48
rect 2203 46 2206 48
rect 2184 43 2191 45
rect 2199 44 2206 46
rect 2184 41 2187 43
rect 2189 41 2191 43
rect 2201 42 2206 44
rect 2208 42 2214 50
rect 2184 36 2191 41
rect 2184 34 2187 36
rect 2189 34 2191 36
rect 2184 32 2191 34
rect 2210 38 2214 42
rect 2267 48 2274 50
rect 2267 46 2269 48
rect 2271 46 2274 48
rect 2267 44 2274 46
rect 2269 42 2274 44
rect 2276 42 2282 50
rect 2245 38 2250 40
rect 2210 34 2216 38
rect 2171 26 2180 32
rect 2171 24 2176 26
rect 2178 24 2180 26
rect 2209 26 2216 34
rect 2171 22 2180 24
rect 2209 24 2211 26
rect 2213 24 2216 26
rect 2209 22 2216 24
rect 2218 22 2223 38
rect 2225 36 2233 38
rect 2225 34 2228 36
rect 2230 34 2233 36
rect 2225 22 2233 34
rect 2235 22 2240 38
rect 2242 26 2250 38
rect 2242 24 2245 26
rect 2247 24 2250 26
rect 2242 22 2250 24
rect 2252 35 2257 40
rect 2278 38 2282 42
rect 2313 38 2318 40
rect 2252 33 2259 35
rect 2278 34 2284 38
rect 2252 31 2255 33
rect 2257 31 2259 33
rect 2252 29 2259 31
rect 2252 22 2257 29
rect 2277 26 2284 34
rect 2277 24 2279 26
rect 2281 24 2284 26
rect 2277 22 2284 24
rect 2286 22 2291 38
rect 2293 36 2301 38
rect 2293 34 2296 36
rect 2298 34 2301 36
rect 2293 22 2301 34
rect 2303 22 2308 38
rect 2310 26 2318 38
rect 2310 24 2313 26
rect 2315 24 2318 26
rect 2310 22 2318 24
rect 2320 35 2325 40
rect 2320 33 2327 35
rect 2320 31 2323 33
rect 2325 31 2327 33
rect 2320 29 2327 31
rect 2320 22 2325 29
rect 8 1 15 3
rect 8 -1 10 1
rect 12 -1 15 1
rect 8 -10 15 -1
rect 17 1 25 3
rect 17 -1 20 1
rect 22 -1 25 1
rect 17 -6 25 -1
rect 17 -8 20 -6
rect 22 -8 25 -6
rect 17 -10 25 -8
rect 27 1 33 3
rect 48 1 55 3
rect 27 -1 35 1
rect 27 -3 30 -1
rect 32 -3 35 -1
rect 27 -10 35 -3
rect 29 -17 35 -10
rect 37 -4 42 1
rect 48 -1 50 1
rect 52 -1 55 1
rect 37 -6 44 -4
rect 37 -8 40 -6
rect 42 -8 44 -6
rect 37 -13 44 -8
rect 48 -10 55 -1
rect 57 1 65 3
rect 57 -1 60 1
rect 62 -1 65 1
rect 57 -6 65 -1
rect 57 -8 60 -6
rect 62 -8 65 -6
rect 57 -10 65 -8
rect 67 1 73 3
rect 67 -1 75 1
rect 67 -3 70 -1
rect 72 -3 75 -1
rect 67 -10 75 -3
rect 37 -15 40 -13
rect 42 -15 44 -13
rect 37 -17 44 -15
rect 69 -17 75 -10
rect 77 -4 82 1
rect 90 -2 95 10
rect 88 -4 95 -2
rect 77 -6 84 -4
rect 77 -8 80 -6
rect 82 -8 84 -6
rect 77 -13 84 -8
rect 77 -15 80 -13
rect 82 -15 84 -13
rect 88 -6 90 -4
rect 92 -6 95 -4
rect 88 -11 95 -6
rect 88 -13 90 -11
rect 92 -13 95 -11
rect 88 -15 95 -13
rect 97 8 106 10
rect 97 6 101 8
rect 103 6 106 8
rect 129 8 143 10
rect 129 7 136 8
rect 97 -2 106 6
rect 113 -2 118 7
rect 97 -15 108 -2
rect 110 -11 118 -2
rect 110 -13 113 -11
rect 115 -13 118 -11
rect 110 -15 118 -13
rect 77 -17 84 -15
rect 113 -18 118 -15
rect 120 -18 125 7
rect 127 6 136 7
rect 138 6 143 8
rect 127 1 143 6
rect 127 -1 136 1
rect 138 -1 143 1
rect 127 -18 143 -1
rect 145 0 153 10
rect 145 -2 148 0
rect 150 -2 153 0
rect 145 -7 153 -2
rect 145 -9 148 -7
rect 150 -9 153 -7
rect 145 -18 153 -9
rect 155 8 163 10
rect 155 6 158 8
rect 160 6 163 8
rect 155 1 163 6
rect 155 -1 158 1
rect 160 -1 163 1
rect 155 -18 163 -1
rect 165 -5 170 10
rect 180 -5 185 10
rect 165 -7 172 -5
rect 165 -9 168 -7
rect 170 -9 172 -7
rect 165 -14 172 -9
rect 165 -16 168 -14
rect 170 -16 172 -14
rect 165 -18 172 -16
rect 178 -7 185 -5
rect 178 -9 180 -7
rect 182 -9 185 -7
rect 178 -14 185 -9
rect 178 -16 180 -14
rect 182 -16 185 -14
rect 178 -18 185 -16
rect 187 8 195 10
rect 187 6 190 8
rect 192 6 195 8
rect 187 1 195 6
rect 187 -1 190 1
rect 192 -1 195 1
rect 187 -18 195 -1
rect 197 0 205 10
rect 197 -2 200 0
rect 202 -2 205 0
rect 197 -7 205 -2
rect 197 -9 200 -7
rect 202 -9 205 -7
rect 197 -18 205 -9
rect 207 8 221 10
rect 207 6 212 8
rect 214 7 221 8
rect 244 8 253 10
rect 214 6 223 7
rect 207 1 223 6
rect 207 -1 212 1
rect 214 -1 223 1
rect 207 -18 223 -1
rect 225 -18 230 7
rect 232 -2 237 7
rect 244 6 247 8
rect 249 6 253 8
rect 244 -2 253 6
rect 232 -11 240 -2
rect 232 -13 235 -11
rect 237 -13 240 -11
rect 232 -15 240 -13
rect 242 -15 253 -2
rect 255 -2 260 10
rect 269 3 274 10
rect 267 1 274 3
rect 267 -1 269 1
rect 271 -1 274 1
rect 255 -4 262 -2
rect 267 -3 274 -1
rect 255 -6 258 -4
rect 260 -6 262 -4
rect 255 -11 262 -6
rect 269 -11 274 -3
rect 276 -11 281 10
rect 283 8 292 10
rect 283 6 288 8
rect 290 6 292 8
rect 283 0 292 6
rect 315 1 322 3
rect 283 -11 294 0
rect 255 -13 258 -11
rect 260 -13 262 -11
rect 255 -15 262 -13
rect 232 -18 237 -15
rect 286 -18 294 -11
rect 296 -2 303 0
rect 296 -4 299 -2
rect 301 -4 303 -2
rect 296 -9 303 -4
rect 296 -11 299 -9
rect 301 -11 303 -9
rect 315 -1 317 1
rect 319 -1 322 1
rect 315 -10 322 -1
rect 324 1 332 3
rect 324 -1 327 1
rect 329 -1 332 1
rect 324 -6 332 -1
rect 324 -8 327 -6
rect 329 -8 332 -6
rect 324 -10 332 -8
rect 334 1 340 3
rect 334 -1 342 1
rect 334 -3 337 -1
rect 339 -3 342 -1
rect 334 -10 342 -3
rect 296 -13 303 -11
rect 296 -18 301 -13
rect 336 -17 342 -10
rect 344 -4 349 1
rect 357 -2 362 10
rect 355 -4 362 -2
rect 344 -6 351 -4
rect 344 -8 347 -6
rect 349 -8 351 -6
rect 344 -13 351 -8
rect 344 -15 347 -13
rect 349 -15 351 -13
rect 355 -6 357 -4
rect 359 -6 362 -4
rect 355 -11 362 -6
rect 355 -13 357 -11
rect 359 -13 362 -11
rect 355 -15 362 -13
rect 364 8 373 10
rect 364 6 368 8
rect 370 6 373 8
rect 396 8 410 10
rect 396 7 403 8
rect 364 -2 373 6
rect 380 -2 385 7
rect 364 -15 375 -2
rect 377 -11 385 -2
rect 377 -13 380 -11
rect 382 -13 385 -11
rect 377 -15 385 -13
rect 344 -17 351 -15
rect 380 -18 385 -15
rect 387 -18 392 7
rect 394 6 403 7
rect 405 6 410 8
rect 394 1 410 6
rect 394 -1 403 1
rect 405 -1 410 1
rect 394 -18 410 -1
rect 412 0 420 10
rect 412 -2 415 0
rect 417 -2 420 0
rect 412 -7 420 -2
rect 412 -9 415 -7
rect 417 -9 420 -7
rect 412 -18 420 -9
rect 422 8 430 10
rect 422 6 425 8
rect 427 6 430 8
rect 422 1 430 6
rect 422 -1 425 1
rect 427 -1 430 1
rect 422 -18 430 -1
rect 432 -5 437 10
rect 447 -5 452 10
rect 432 -7 439 -5
rect 432 -9 435 -7
rect 437 -9 439 -7
rect 432 -14 439 -9
rect 432 -16 435 -14
rect 437 -16 439 -14
rect 432 -18 439 -16
rect 445 -7 452 -5
rect 445 -9 447 -7
rect 449 -9 452 -7
rect 445 -14 452 -9
rect 445 -16 447 -14
rect 449 -16 452 -14
rect 445 -18 452 -16
rect 454 8 462 10
rect 454 6 457 8
rect 459 6 462 8
rect 454 1 462 6
rect 454 -1 457 1
rect 459 -1 462 1
rect 454 -18 462 -1
rect 464 0 472 10
rect 464 -2 467 0
rect 469 -2 472 0
rect 464 -7 472 -2
rect 464 -9 467 -7
rect 469 -9 472 -7
rect 464 -18 472 -9
rect 474 8 488 10
rect 474 6 479 8
rect 481 7 488 8
rect 511 8 520 10
rect 481 6 490 7
rect 474 1 490 6
rect 474 -1 479 1
rect 481 -1 490 1
rect 474 -18 490 -1
rect 492 -18 497 7
rect 499 -2 504 7
rect 511 6 514 8
rect 516 6 520 8
rect 511 -2 520 6
rect 499 -11 507 -2
rect 499 -13 502 -11
rect 504 -13 507 -11
rect 499 -15 507 -13
rect 509 -15 520 -2
rect 522 -2 527 10
rect 536 3 541 10
rect 534 1 541 3
rect 534 -1 536 1
rect 538 -1 541 1
rect 522 -4 529 -2
rect 534 -3 541 -1
rect 522 -6 525 -4
rect 527 -6 529 -4
rect 522 -11 529 -6
rect 536 -11 541 -3
rect 543 -11 548 10
rect 550 8 559 10
rect 550 6 555 8
rect 557 6 559 8
rect 550 0 559 6
rect 582 1 589 3
rect 550 -11 561 0
rect 522 -13 525 -11
rect 527 -13 529 -11
rect 522 -15 529 -13
rect 499 -18 504 -15
rect 553 -18 561 -11
rect 563 -2 570 0
rect 563 -4 566 -2
rect 568 -4 570 -2
rect 563 -9 570 -4
rect 563 -11 566 -9
rect 568 -11 570 -9
rect 582 -1 584 1
rect 586 -1 589 1
rect 582 -10 589 -1
rect 591 1 599 3
rect 591 -1 594 1
rect 596 -1 599 1
rect 591 -6 599 -1
rect 591 -8 594 -6
rect 596 -8 599 -6
rect 591 -10 599 -8
rect 601 1 607 3
rect 601 -1 609 1
rect 601 -3 604 -1
rect 606 -3 609 -1
rect 601 -10 609 -3
rect 563 -13 570 -11
rect 563 -18 568 -13
rect 603 -17 609 -10
rect 611 -4 616 1
rect 624 -2 629 10
rect 622 -4 629 -2
rect 611 -6 618 -4
rect 611 -8 614 -6
rect 616 -8 618 -6
rect 611 -13 618 -8
rect 611 -15 614 -13
rect 616 -15 618 -13
rect 622 -6 624 -4
rect 626 -6 629 -4
rect 622 -11 629 -6
rect 622 -13 624 -11
rect 626 -13 629 -11
rect 622 -15 629 -13
rect 631 8 640 10
rect 631 6 635 8
rect 637 6 640 8
rect 663 8 677 10
rect 663 7 670 8
rect 631 -2 640 6
rect 647 -2 652 7
rect 631 -15 642 -2
rect 644 -11 652 -2
rect 644 -13 647 -11
rect 649 -13 652 -11
rect 644 -15 652 -13
rect 611 -17 618 -15
rect 647 -18 652 -15
rect 654 -18 659 7
rect 661 6 670 7
rect 672 6 677 8
rect 661 1 677 6
rect 661 -1 670 1
rect 672 -1 677 1
rect 661 -18 677 -1
rect 679 0 687 10
rect 679 -2 682 0
rect 684 -2 687 0
rect 679 -7 687 -2
rect 679 -9 682 -7
rect 684 -9 687 -7
rect 679 -18 687 -9
rect 689 8 697 10
rect 689 6 692 8
rect 694 6 697 8
rect 689 1 697 6
rect 689 -1 692 1
rect 694 -1 697 1
rect 689 -18 697 -1
rect 699 -5 704 10
rect 714 -5 719 10
rect 699 -7 706 -5
rect 699 -9 702 -7
rect 704 -9 706 -7
rect 699 -14 706 -9
rect 699 -16 702 -14
rect 704 -16 706 -14
rect 699 -18 706 -16
rect 712 -7 719 -5
rect 712 -9 714 -7
rect 716 -9 719 -7
rect 712 -14 719 -9
rect 712 -16 714 -14
rect 716 -16 719 -14
rect 712 -18 719 -16
rect 721 8 729 10
rect 721 6 724 8
rect 726 6 729 8
rect 721 1 729 6
rect 721 -1 724 1
rect 726 -1 729 1
rect 721 -18 729 -1
rect 731 0 739 10
rect 731 -2 734 0
rect 736 -2 739 0
rect 731 -7 739 -2
rect 731 -9 734 -7
rect 736 -9 739 -7
rect 731 -18 739 -9
rect 741 8 755 10
rect 741 6 746 8
rect 748 7 755 8
rect 778 8 787 10
rect 748 6 757 7
rect 741 1 757 6
rect 741 -1 746 1
rect 748 -1 757 1
rect 741 -18 757 -1
rect 759 -18 764 7
rect 766 -2 771 7
rect 778 6 781 8
rect 783 6 787 8
rect 778 -2 787 6
rect 766 -11 774 -2
rect 766 -13 769 -11
rect 771 -13 774 -11
rect 766 -15 774 -13
rect 776 -15 787 -2
rect 789 -2 794 10
rect 803 3 808 10
rect 801 1 808 3
rect 801 -1 803 1
rect 805 -1 808 1
rect 789 -4 796 -2
rect 801 -3 808 -1
rect 789 -6 792 -4
rect 794 -6 796 -4
rect 789 -11 796 -6
rect 803 -11 808 -3
rect 810 -11 815 10
rect 817 8 826 10
rect 817 6 822 8
rect 824 6 826 8
rect 817 0 826 6
rect 849 1 856 3
rect 817 -11 828 0
rect 789 -13 792 -11
rect 794 -13 796 -11
rect 789 -15 796 -13
rect 766 -18 771 -15
rect 820 -18 828 -11
rect 830 -2 837 0
rect 830 -4 833 -2
rect 835 -4 837 -2
rect 830 -9 837 -4
rect 830 -11 833 -9
rect 835 -11 837 -9
rect 849 -1 851 1
rect 853 -1 856 1
rect 849 -10 856 -1
rect 858 1 866 3
rect 858 -1 861 1
rect 863 -1 866 1
rect 858 -6 866 -1
rect 858 -8 861 -6
rect 863 -8 866 -6
rect 858 -10 866 -8
rect 868 1 874 3
rect 868 -1 876 1
rect 868 -3 871 -1
rect 873 -3 876 -1
rect 868 -10 876 -3
rect 830 -13 837 -11
rect 830 -18 835 -13
rect 870 -17 876 -10
rect 878 -4 883 1
rect 891 -2 896 10
rect 889 -4 896 -2
rect 878 -6 885 -4
rect 878 -8 881 -6
rect 883 -8 885 -6
rect 878 -13 885 -8
rect 878 -15 881 -13
rect 883 -15 885 -13
rect 889 -6 891 -4
rect 893 -6 896 -4
rect 889 -11 896 -6
rect 889 -13 891 -11
rect 893 -13 896 -11
rect 889 -15 896 -13
rect 898 8 907 10
rect 898 6 902 8
rect 904 6 907 8
rect 930 8 944 10
rect 930 7 937 8
rect 898 -2 907 6
rect 914 -2 919 7
rect 898 -15 909 -2
rect 911 -11 919 -2
rect 911 -13 914 -11
rect 916 -13 919 -11
rect 911 -15 919 -13
rect 878 -17 885 -15
rect 914 -18 919 -15
rect 921 -18 926 7
rect 928 6 937 7
rect 939 6 944 8
rect 928 1 944 6
rect 928 -1 937 1
rect 939 -1 944 1
rect 928 -18 944 -1
rect 946 0 954 10
rect 946 -2 949 0
rect 951 -2 954 0
rect 946 -7 954 -2
rect 946 -9 949 -7
rect 951 -9 954 -7
rect 946 -18 954 -9
rect 956 8 964 10
rect 956 6 959 8
rect 961 6 964 8
rect 956 1 964 6
rect 956 -1 959 1
rect 961 -1 964 1
rect 956 -18 964 -1
rect 966 -5 971 10
rect 981 -5 986 10
rect 966 -7 973 -5
rect 966 -9 969 -7
rect 971 -9 973 -7
rect 966 -14 973 -9
rect 966 -16 969 -14
rect 971 -16 973 -14
rect 966 -18 973 -16
rect 979 -7 986 -5
rect 979 -9 981 -7
rect 983 -9 986 -7
rect 979 -14 986 -9
rect 979 -16 981 -14
rect 983 -16 986 -14
rect 979 -18 986 -16
rect 988 8 996 10
rect 988 6 991 8
rect 993 6 996 8
rect 988 1 996 6
rect 988 -1 991 1
rect 993 -1 996 1
rect 988 -18 996 -1
rect 998 0 1006 10
rect 998 -2 1001 0
rect 1003 -2 1006 0
rect 998 -7 1006 -2
rect 998 -9 1001 -7
rect 1003 -9 1006 -7
rect 998 -18 1006 -9
rect 1008 8 1022 10
rect 1008 6 1013 8
rect 1015 7 1022 8
rect 1045 8 1054 10
rect 1015 6 1024 7
rect 1008 1 1024 6
rect 1008 -1 1013 1
rect 1015 -1 1024 1
rect 1008 -18 1024 -1
rect 1026 -18 1031 7
rect 1033 -2 1038 7
rect 1045 6 1048 8
rect 1050 6 1054 8
rect 1045 -2 1054 6
rect 1033 -11 1041 -2
rect 1033 -13 1036 -11
rect 1038 -13 1041 -11
rect 1033 -15 1041 -13
rect 1043 -15 1054 -2
rect 1056 -2 1061 10
rect 1070 3 1075 10
rect 1068 1 1075 3
rect 1068 -1 1070 1
rect 1072 -1 1075 1
rect 1056 -4 1063 -2
rect 1068 -3 1075 -1
rect 1056 -6 1059 -4
rect 1061 -6 1063 -4
rect 1056 -11 1063 -6
rect 1070 -11 1075 -3
rect 1077 -11 1082 10
rect 1084 8 1093 10
rect 1084 6 1089 8
rect 1091 6 1093 8
rect 1084 0 1093 6
rect 1116 1 1123 3
rect 1084 -11 1095 0
rect 1056 -13 1059 -11
rect 1061 -13 1063 -11
rect 1056 -15 1063 -13
rect 1033 -18 1038 -15
rect 1087 -18 1095 -11
rect 1097 -2 1104 0
rect 1097 -4 1100 -2
rect 1102 -4 1104 -2
rect 1097 -9 1104 -4
rect 1097 -11 1100 -9
rect 1102 -11 1104 -9
rect 1116 -1 1118 1
rect 1120 -1 1123 1
rect 1116 -10 1123 -1
rect 1125 1 1133 3
rect 1125 -1 1128 1
rect 1130 -1 1133 1
rect 1125 -6 1133 -1
rect 1125 -8 1128 -6
rect 1130 -8 1133 -6
rect 1125 -10 1133 -8
rect 1135 1 1141 3
rect 1135 -1 1143 1
rect 1135 -3 1138 -1
rect 1140 -3 1143 -1
rect 1135 -10 1143 -3
rect 1097 -13 1104 -11
rect 1097 -18 1102 -13
rect 1137 -17 1143 -10
rect 1145 -4 1150 1
rect 1158 -2 1163 10
rect 1156 -4 1163 -2
rect 1145 -6 1152 -4
rect 1145 -8 1148 -6
rect 1150 -8 1152 -6
rect 1145 -13 1152 -8
rect 1145 -15 1148 -13
rect 1150 -15 1152 -13
rect 1156 -6 1158 -4
rect 1160 -6 1163 -4
rect 1156 -11 1163 -6
rect 1156 -13 1158 -11
rect 1160 -13 1163 -11
rect 1156 -15 1163 -13
rect 1165 8 1174 10
rect 1165 6 1169 8
rect 1171 6 1174 8
rect 1197 8 1211 10
rect 1197 7 1204 8
rect 1165 -2 1174 6
rect 1181 -2 1186 7
rect 1165 -15 1176 -2
rect 1178 -11 1186 -2
rect 1178 -13 1181 -11
rect 1183 -13 1186 -11
rect 1178 -15 1186 -13
rect 1145 -17 1152 -15
rect 1181 -18 1186 -15
rect 1188 -18 1193 7
rect 1195 6 1204 7
rect 1206 6 1211 8
rect 1195 1 1211 6
rect 1195 -1 1204 1
rect 1206 -1 1211 1
rect 1195 -18 1211 -1
rect 1213 0 1221 10
rect 1213 -2 1216 0
rect 1218 -2 1221 0
rect 1213 -7 1221 -2
rect 1213 -9 1216 -7
rect 1218 -9 1221 -7
rect 1213 -18 1221 -9
rect 1223 8 1231 10
rect 1223 6 1226 8
rect 1228 6 1231 8
rect 1223 1 1231 6
rect 1223 -1 1226 1
rect 1228 -1 1231 1
rect 1223 -18 1231 -1
rect 1233 -5 1238 10
rect 1248 -5 1253 10
rect 1233 -7 1240 -5
rect 1233 -9 1236 -7
rect 1238 -9 1240 -7
rect 1233 -14 1240 -9
rect 1233 -16 1236 -14
rect 1238 -16 1240 -14
rect 1233 -18 1240 -16
rect 1246 -7 1253 -5
rect 1246 -9 1248 -7
rect 1250 -9 1253 -7
rect 1246 -14 1253 -9
rect 1246 -16 1248 -14
rect 1250 -16 1253 -14
rect 1246 -18 1253 -16
rect 1255 8 1263 10
rect 1255 6 1258 8
rect 1260 6 1263 8
rect 1255 1 1263 6
rect 1255 -1 1258 1
rect 1260 -1 1263 1
rect 1255 -18 1263 -1
rect 1265 0 1273 10
rect 1265 -2 1268 0
rect 1270 -2 1273 0
rect 1265 -7 1273 -2
rect 1265 -9 1268 -7
rect 1270 -9 1273 -7
rect 1265 -18 1273 -9
rect 1275 8 1289 10
rect 1275 6 1280 8
rect 1282 7 1289 8
rect 1312 8 1321 10
rect 1282 6 1291 7
rect 1275 1 1291 6
rect 1275 -1 1280 1
rect 1282 -1 1291 1
rect 1275 -18 1291 -1
rect 1293 -18 1298 7
rect 1300 -2 1305 7
rect 1312 6 1315 8
rect 1317 6 1321 8
rect 1312 -2 1321 6
rect 1300 -11 1308 -2
rect 1300 -13 1303 -11
rect 1305 -13 1308 -11
rect 1300 -15 1308 -13
rect 1310 -15 1321 -2
rect 1323 -2 1328 10
rect 1337 3 1342 10
rect 1335 1 1342 3
rect 1335 -1 1337 1
rect 1339 -1 1342 1
rect 1323 -4 1330 -2
rect 1335 -3 1342 -1
rect 1323 -6 1326 -4
rect 1328 -6 1330 -4
rect 1323 -11 1330 -6
rect 1337 -11 1342 -3
rect 1344 -11 1349 10
rect 1351 8 1360 10
rect 1351 6 1356 8
rect 1358 6 1360 8
rect 1351 0 1360 6
rect 1383 1 1390 3
rect 1351 -11 1362 0
rect 1323 -13 1326 -11
rect 1328 -13 1330 -11
rect 1323 -15 1330 -13
rect 1300 -18 1305 -15
rect 1354 -18 1362 -11
rect 1364 -2 1371 0
rect 1364 -4 1367 -2
rect 1369 -4 1371 -2
rect 1364 -9 1371 -4
rect 1364 -11 1367 -9
rect 1369 -11 1371 -9
rect 1383 -1 1385 1
rect 1387 -1 1390 1
rect 1383 -10 1390 -1
rect 1392 1 1400 3
rect 1392 -1 1395 1
rect 1397 -1 1400 1
rect 1392 -6 1400 -1
rect 1392 -8 1395 -6
rect 1397 -8 1400 -6
rect 1392 -10 1400 -8
rect 1402 1 1408 3
rect 1402 -1 1410 1
rect 1402 -3 1405 -1
rect 1407 -3 1410 -1
rect 1402 -10 1410 -3
rect 1364 -13 1371 -11
rect 1364 -18 1369 -13
rect 1404 -17 1410 -10
rect 1412 -4 1417 1
rect 1425 -2 1430 10
rect 1423 -4 1430 -2
rect 1412 -6 1419 -4
rect 1412 -8 1415 -6
rect 1417 -8 1419 -6
rect 1412 -13 1419 -8
rect 1412 -15 1415 -13
rect 1417 -15 1419 -13
rect 1423 -6 1425 -4
rect 1427 -6 1430 -4
rect 1423 -11 1430 -6
rect 1423 -13 1425 -11
rect 1427 -13 1430 -11
rect 1423 -15 1430 -13
rect 1432 8 1441 10
rect 1432 6 1436 8
rect 1438 6 1441 8
rect 1464 8 1478 10
rect 1464 7 1471 8
rect 1432 -2 1441 6
rect 1448 -2 1453 7
rect 1432 -15 1443 -2
rect 1445 -11 1453 -2
rect 1445 -13 1448 -11
rect 1450 -13 1453 -11
rect 1445 -15 1453 -13
rect 1412 -17 1419 -15
rect 1448 -18 1453 -15
rect 1455 -18 1460 7
rect 1462 6 1471 7
rect 1473 6 1478 8
rect 1462 1 1478 6
rect 1462 -1 1471 1
rect 1473 -1 1478 1
rect 1462 -18 1478 -1
rect 1480 0 1488 10
rect 1480 -2 1483 0
rect 1485 -2 1488 0
rect 1480 -7 1488 -2
rect 1480 -9 1483 -7
rect 1485 -9 1488 -7
rect 1480 -18 1488 -9
rect 1490 8 1498 10
rect 1490 6 1493 8
rect 1495 6 1498 8
rect 1490 1 1498 6
rect 1490 -1 1493 1
rect 1495 -1 1498 1
rect 1490 -18 1498 -1
rect 1500 -5 1505 10
rect 1515 -5 1520 10
rect 1500 -7 1507 -5
rect 1500 -9 1503 -7
rect 1505 -9 1507 -7
rect 1500 -14 1507 -9
rect 1500 -16 1503 -14
rect 1505 -16 1507 -14
rect 1500 -18 1507 -16
rect 1513 -7 1520 -5
rect 1513 -9 1515 -7
rect 1517 -9 1520 -7
rect 1513 -14 1520 -9
rect 1513 -16 1515 -14
rect 1517 -16 1520 -14
rect 1513 -18 1520 -16
rect 1522 8 1530 10
rect 1522 6 1525 8
rect 1527 6 1530 8
rect 1522 1 1530 6
rect 1522 -1 1525 1
rect 1527 -1 1530 1
rect 1522 -18 1530 -1
rect 1532 0 1540 10
rect 1532 -2 1535 0
rect 1537 -2 1540 0
rect 1532 -7 1540 -2
rect 1532 -9 1535 -7
rect 1537 -9 1540 -7
rect 1532 -18 1540 -9
rect 1542 8 1556 10
rect 1542 6 1547 8
rect 1549 7 1556 8
rect 1579 8 1588 10
rect 1549 6 1558 7
rect 1542 1 1558 6
rect 1542 -1 1547 1
rect 1549 -1 1558 1
rect 1542 -18 1558 -1
rect 1560 -18 1565 7
rect 1567 -2 1572 7
rect 1579 6 1582 8
rect 1584 6 1588 8
rect 1579 -2 1588 6
rect 1567 -11 1575 -2
rect 1567 -13 1570 -11
rect 1572 -13 1575 -11
rect 1567 -15 1575 -13
rect 1577 -15 1588 -2
rect 1590 -2 1595 10
rect 1604 3 1609 10
rect 1602 1 1609 3
rect 1602 -1 1604 1
rect 1606 -1 1609 1
rect 1590 -4 1597 -2
rect 1602 -3 1609 -1
rect 1590 -6 1593 -4
rect 1595 -6 1597 -4
rect 1590 -11 1597 -6
rect 1604 -11 1609 -3
rect 1611 -11 1616 10
rect 1618 8 1627 10
rect 1618 6 1623 8
rect 1625 6 1627 8
rect 1618 0 1627 6
rect 1650 1 1657 3
rect 1618 -11 1629 0
rect 1590 -13 1593 -11
rect 1595 -13 1597 -11
rect 1590 -15 1597 -13
rect 1567 -18 1572 -15
rect 1621 -18 1629 -11
rect 1631 -2 1638 0
rect 1631 -4 1634 -2
rect 1636 -4 1638 -2
rect 1631 -9 1638 -4
rect 1631 -11 1634 -9
rect 1636 -11 1638 -9
rect 1650 -1 1652 1
rect 1654 -1 1657 1
rect 1650 -10 1657 -1
rect 1659 1 1667 3
rect 1659 -1 1662 1
rect 1664 -1 1667 1
rect 1659 -6 1667 -1
rect 1659 -8 1662 -6
rect 1664 -8 1667 -6
rect 1659 -10 1667 -8
rect 1669 1 1675 3
rect 1669 -1 1677 1
rect 1669 -3 1672 -1
rect 1674 -3 1677 -1
rect 1669 -10 1677 -3
rect 1631 -13 1638 -11
rect 1631 -18 1636 -13
rect 1671 -17 1677 -10
rect 1679 -4 1684 1
rect 1692 -2 1697 10
rect 1690 -4 1697 -2
rect 1679 -6 1686 -4
rect 1679 -8 1682 -6
rect 1684 -8 1686 -6
rect 1679 -13 1686 -8
rect 1679 -15 1682 -13
rect 1684 -15 1686 -13
rect 1690 -6 1692 -4
rect 1694 -6 1697 -4
rect 1690 -11 1697 -6
rect 1690 -13 1692 -11
rect 1694 -13 1697 -11
rect 1690 -15 1697 -13
rect 1699 8 1708 10
rect 1699 6 1703 8
rect 1705 6 1708 8
rect 1731 8 1745 10
rect 1731 7 1738 8
rect 1699 -2 1708 6
rect 1715 -2 1720 7
rect 1699 -15 1710 -2
rect 1712 -11 1720 -2
rect 1712 -13 1715 -11
rect 1717 -13 1720 -11
rect 1712 -15 1720 -13
rect 1679 -17 1686 -15
rect 1715 -18 1720 -15
rect 1722 -18 1727 7
rect 1729 6 1738 7
rect 1740 6 1745 8
rect 1729 1 1745 6
rect 1729 -1 1738 1
rect 1740 -1 1745 1
rect 1729 -18 1745 -1
rect 1747 0 1755 10
rect 1747 -2 1750 0
rect 1752 -2 1755 0
rect 1747 -7 1755 -2
rect 1747 -9 1750 -7
rect 1752 -9 1755 -7
rect 1747 -18 1755 -9
rect 1757 8 1765 10
rect 1757 6 1760 8
rect 1762 6 1765 8
rect 1757 1 1765 6
rect 1757 -1 1760 1
rect 1762 -1 1765 1
rect 1757 -18 1765 -1
rect 1767 -5 1772 10
rect 1782 -5 1787 10
rect 1767 -7 1774 -5
rect 1767 -9 1770 -7
rect 1772 -9 1774 -7
rect 1767 -14 1774 -9
rect 1767 -16 1770 -14
rect 1772 -16 1774 -14
rect 1767 -18 1774 -16
rect 1780 -7 1787 -5
rect 1780 -9 1782 -7
rect 1784 -9 1787 -7
rect 1780 -14 1787 -9
rect 1780 -16 1782 -14
rect 1784 -16 1787 -14
rect 1780 -18 1787 -16
rect 1789 8 1797 10
rect 1789 6 1792 8
rect 1794 6 1797 8
rect 1789 1 1797 6
rect 1789 -1 1792 1
rect 1794 -1 1797 1
rect 1789 -18 1797 -1
rect 1799 0 1807 10
rect 1799 -2 1802 0
rect 1804 -2 1807 0
rect 1799 -7 1807 -2
rect 1799 -9 1802 -7
rect 1804 -9 1807 -7
rect 1799 -18 1807 -9
rect 1809 8 1823 10
rect 1809 6 1814 8
rect 1816 7 1823 8
rect 1846 8 1855 10
rect 1816 6 1825 7
rect 1809 1 1825 6
rect 1809 -1 1814 1
rect 1816 -1 1825 1
rect 1809 -18 1825 -1
rect 1827 -18 1832 7
rect 1834 -2 1839 7
rect 1846 6 1849 8
rect 1851 6 1855 8
rect 1846 -2 1855 6
rect 1834 -11 1842 -2
rect 1834 -13 1837 -11
rect 1839 -13 1842 -11
rect 1834 -15 1842 -13
rect 1844 -15 1855 -2
rect 1857 -2 1862 10
rect 1871 3 1876 10
rect 1869 1 1876 3
rect 1869 -1 1871 1
rect 1873 -1 1876 1
rect 1857 -4 1864 -2
rect 1869 -3 1876 -1
rect 1857 -6 1860 -4
rect 1862 -6 1864 -4
rect 1857 -11 1864 -6
rect 1871 -11 1876 -3
rect 1878 -11 1883 10
rect 1885 8 1894 10
rect 1885 6 1890 8
rect 1892 6 1894 8
rect 1885 0 1894 6
rect 1885 -11 1896 0
rect 1857 -13 1860 -11
rect 1862 -13 1864 -11
rect 1857 -15 1864 -13
rect 1834 -18 1839 -15
rect 1888 -18 1896 -11
rect 1898 -2 1905 0
rect 1898 -4 1901 -2
rect 1903 -4 1905 -2
rect 1898 -9 1905 -4
rect 1898 -11 1901 -9
rect 1903 -11 1905 -9
rect 1922 -11 1927 10
rect 1898 -13 1905 -11
rect 1920 -13 1927 -11
rect 1898 -18 1903 -13
rect 1920 -15 1922 -13
rect 1924 -15 1927 -13
rect 1920 -17 1927 -15
rect 1929 8 1941 10
rect 1929 6 1932 8
rect 1934 6 1941 8
rect 1929 1 1941 6
rect 1958 1 1963 10
rect 1929 -1 1932 1
rect 1934 -1 1943 1
rect 1929 -17 1943 -1
rect 1945 -6 1953 1
rect 1945 -8 1948 -6
rect 1950 -8 1953 -6
rect 1945 -13 1953 -8
rect 1945 -15 1948 -13
rect 1950 -15 1953 -13
rect 1945 -17 1953 -15
rect 1955 -6 1963 1
rect 1955 -8 1958 -6
rect 1960 -8 1963 -6
rect 1955 -17 1963 -8
rect 1965 4 1970 10
rect 1965 2 1972 4
rect 1965 0 1968 2
rect 1970 0 1972 2
rect 1965 -2 1972 0
rect 1978 -2 1983 10
rect 1965 -17 1970 -2
rect 1976 -4 1983 -2
rect 1976 -6 1978 -4
rect 1980 -6 1983 -4
rect 1976 -11 1983 -6
rect 1976 -13 1978 -11
rect 1980 -13 1983 -11
rect 1976 -15 1983 -13
rect 1985 8 1994 10
rect 1985 6 1989 8
rect 1991 6 1994 8
rect 2017 8 2031 10
rect 2017 7 2024 8
rect 1985 -2 1994 6
rect 2001 -2 2006 7
rect 1985 -15 1996 -2
rect 1998 -11 2006 -2
rect 1998 -13 2001 -11
rect 2003 -13 2006 -11
rect 1998 -15 2006 -13
rect 2001 -18 2006 -15
rect 2008 -18 2013 7
rect 2015 6 2024 7
rect 2026 6 2031 8
rect 2015 1 2031 6
rect 2015 -1 2024 1
rect 2026 -1 2031 1
rect 2015 -18 2031 -1
rect 2033 0 2041 10
rect 2033 -2 2036 0
rect 2038 -2 2041 0
rect 2033 -7 2041 -2
rect 2033 -9 2036 -7
rect 2038 -9 2041 -7
rect 2033 -18 2041 -9
rect 2043 8 2051 10
rect 2043 6 2046 8
rect 2048 6 2051 8
rect 2043 1 2051 6
rect 2043 -1 2046 1
rect 2048 -1 2051 1
rect 2043 -18 2051 -1
rect 2053 -5 2058 10
rect 2068 -5 2073 10
rect 2053 -7 2060 -5
rect 2053 -9 2056 -7
rect 2058 -9 2060 -7
rect 2053 -14 2060 -9
rect 2053 -16 2056 -14
rect 2058 -16 2060 -14
rect 2053 -18 2060 -16
rect 2066 -7 2073 -5
rect 2066 -9 2068 -7
rect 2070 -9 2073 -7
rect 2066 -14 2073 -9
rect 2066 -16 2068 -14
rect 2070 -16 2073 -14
rect 2066 -18 2073 -16
rect 2075 8 2083 10
rect 2075 6 2078 8
rect 2080 6 2083 8
rect 2075 1 2083 6
rect 2075 -1 2078 1
rect 2080 -1 2083 1
rect 2075 -18 2083 -1
rect 2085 0 2093 10
rect 2085 -2 2088 0
rect 2090 -2 2093 0
rect 2085 -7 2093 -2
rect 2085 -9 2088 -7
rect 2090 -9 2093 -7
rect 2085 -18 2093 -9
rect 2095 8 2109 10
rect 2095 6 2100 8
rect 2102 7 2109 8
rect 2132 8 2141 10
rect 2102 6 2111 7
rect 2095 1 2111 6
rect 2095 -1 2100 1
rect 2102 -1 2111 1
rect 2095 -18 2111 -1
rect 2113 -18 2118 7
rect 2120 -2 2125 7
rect 2132 6 2135 8
rect 2137 6 2141 8
rect 2132 -2 2141 6
rect 2120 -11 2128 -2
rect 2120 -13 2123 -11
rect 2125 -13 2128 -11
rect 2120 -15 2128 -13
rect 2130 -15 2141 -2
rect 2143 -2 2148 10
rect 2157 3 2162 10
rect 2155 1 2162 3
rect 2155 -1 2157 1
rect 2159 -1 2162 1
rect 2143 -4 2150 -2
rect 2155 -3 2162 -1
rect 2143 -6 2146 -4
rect 2148 -6 2150 -4
rect 2143 -11 2150 -6
rect 2157 -11 2162 -3
rect 2164 -11 2169 10
rect 2171 8 2180 10
rect 2171 6 2176 8
rect 2178 6 2180 8
rect 2209 8 2216 10
rect 2171 0 2180 6
rect 2209 6 2211 8
rect 2213 6 2216 8
rect 2171 -11 2182 0
rect 2143 -13 2146 -11
rect 2148 -13 2150 -11
rect 2143 -15 2150 -13
rect 2120 -18 2125 -15
rect 2174 -18 2182 -11
rect 2184 -2 2191 0
rect 2184 -4 2187 -2
rect 2189 -4 2191 -2
rect 2184 -9 2191 -4
rect 2209 -2 2216 6
rect 2184 -11 2187 -9
rect 2189 -11 2191 -9
rect 2210 -6 2216 -2
rect 2218 -6 2223 10
rect 2225 -2 2233 10
rect 2225 -4 2228 -2
rect 2230 -4 2233 -2
rect 2225 -6 2233 -4
rect 2235 -6 2240 10
rect 2242 8 2250 10
rect 2242 6 2245 8
rect 2247 6 2250 8
rect 2242 -6 2250 6
rect 2210 -10 2214 -6
rect 2184 -13 2191 -11
rect 2201 -12 2206 -10
rect 2184 -18 2189 -13
rect 2199 -14 2206 -12
rect 2199 -16 2201 -14
rect 2203 -16 2206 -14
rect 2199 -18 2206 -16
rect 2208 -18 2214 -10
rect 2245 -8 2250 -6
rect 2252 3 2257 10
rect 2277 8 2284 10
rect 2277 6 2279 8
rect 2281 6 2284 8
rect 2252 1 2259 3
rect 2252 -1 2255 1
rect 2257 -1 2259 1
rect 2252 -3 2259 -1
rect 2277 -2 2284 6
rect 2252 -8 2257 -3
rect 2278 -6 2284 -2
rect 2286 -6 2291 10
rect 2293 -2 2301 10
rect 2293 -4 2296 -2
rect 2298 -4 2301 -2
rect 2293 -6 2301 -4
rect 2303 -6 2308 10
rect 2310 8 2318 10
rect 2310 6 2313 8
rect 2315 6 2318 8
rect 2310 -6 2318 6
rect 2278 -10 2282 -6
rect 2269 -12 2274 -10
rect 2267 -14 2274 -12
rect 2267 -16 2269 -14
rect 2271 -16 2274 -14
rect 2267 -18 2274 -16
rect 2276 -18 2282 -10
rect 2313 -8 2318 -6
rect 2320 3 2325 10
rect 2320 1 2327 3
rect 2320 -1 2323 1
rect 2325 -1 2327 1
rect 2320 -3 2327 -1
rect 2320 -8 2325 -3
rect 29 -102 35 -95
rect 8 -111 15 -102
rect 8 -113 10 -111
rect 12 -113 15 -111
rect 8 -115 15 -113
rect 17 -104 25 -102
rect 17 -106 20 -104
rect 22 -106 25 -104
rect 17 -111 25 -106
rect 17 -113 20 -111
rect 22 -113 25 -111
rect 17 -115 25 -113
rect 27 -109 35 -102
rect 27 -111 30 -109
rect 32 -111 35 -109
rect 27 -113 35 -111
rect 37 -98 44 -95
rect 37 -100 40 -98
rect 42 -100 44 -98
rect 37 -106 44 -100
rect 69 -102 75 -95
rect 37 -108 40 -106
rect 42 -108 44 -106
rect 37 -110 44 -108
rect 37 -113 42 -110
rect 48 -111 55 -102
rect 48 -113 50 -111
rect 52 -113 55 -111
rect 27 -115 33 -113
rect 48 -115 55 -113
rect 57 -104 65 -102
rect 57 -106 60 -104
rect 62 -106 65 -104
rect 57 -111 65 -106
rect 57 -113 60 -111
rect 62 -113 65 -111
rect 57 -115 65 -113
rect 67 -109 75 -102
rect 67 -111 70 -109
rect 72 -111 75 -109
rect 67 -113 75 -111
rect 77 -97 84 -95
rect 113 -97 118 -94
rect 77 -99 80 -97
rect 82 -99 84 -97
rect 77 -104 84 -99
rect 77 -106 80 -104
rect 82 -106 84 -104
rect 77 -108 84 -106
rect 88 -99 95 -97
rect 88 -101 90 -99
rect 92 -101 95 -99
rect 88 -106 95 -101
rect 88 -108 90 -106
rect 92 -108 95 -106
rect 77 -113 82 -108
rect 88 -110 95 -108
rect 67 -115 73 -113
rect 90 -122 95 -110
rect 97 -110 108 -97
rect 110 -99 118 -97
rect 110 -101 113 -99
rect 115 -101 118 -99
rect 110 -110 118 -101
rect 97 -118 106 -110
rect 97 -120 101 -118
rect 103 -120 106 -118
rect 113 -119 118 -110
rect 120 -119 125 -94
rect 127 -111 143 -94
rect 127 -113 136 -111
rect 138 -113 143 -111
rect 127 -118 143 -113
rect 127 -119 136 -118
rect 97 -122 106 -120
rect 129 -120 136 -119
rect 138 -120 143 -118
rect 129 -122 143 -120
rect 145 -103 153 -94
rect 145 -105 148 -103
rect 150 -105 153 -103
rect 145 -110 153 -105
rect 145 -112 148 -110
rect 150 -112 153 -110
rect 145 -122 153 -112
rect 155 -111 163 -94
rect 155 -113 158 -111
rect 160 -113 163 -111
rect 155 -118 163 -113
rect 155 -120 158 -118
rect 160 -120 163 -118
rect 155 -122 163 -120
rect 165 -96 172 -94
rect 165 -98 168 -96
rect 170 -98 172 -96
rect 165 -103 172 -98
rect 165 -105 168 -103
rect 170 -105 172 -103
rect 165 -107 172 -105
rect 178 -96 185 -94
rect 178 -98 180 -96
rect 182 -98 185 -96
rect 178 -103 185 -98
rect 178 -105 180 -103
rect 182 -105 185 -103
rect 178 -107 185 -105
rect 165 -122 170 -107
rect 180 -122 185 -107
rect 187 -111 195 -94
rect 187 -113 190 -111
rect 192 -113 195 -111
rect 187 -118 195 -113
rect 187 -120 190 -118
rect 192 -120 195 -118
rect 187 -122 195 -120
rect 197 -103 205 -94
rect 197 -105 200 -103
rect 202 -105 205 -103
rect 197 -110 205 -105
rect 197 -112 200 -110
rect 202 -112 205 -110
rect 197 -122 205 -112
rect 207 -111 223 -94
rect 207 -113 212 -111
rect 214 -113 223 -111
rect 207 -118 223 -113
rect 207 -120 212 -118
rect 214 -119 223 -118
rect 225 -119 230 -94
rect 232 -97 237 -94
rect 232 -99 240 -97
rect 232 -101 235 -99
rect 237 -101 240 -99
rect 232 -110 240 -101
rect 242 -110 253 -97
rect 232 -119 237 -110
rect 244 -118 253 -110
rect 214 -120 221 -119
rect 207 -122 221 -120
rect 244 -120 247 -118
rect 249 -120 253 -118
rect 244 -122 253 -120
rect 255 -99 262 -97
rect 255 -101 258 -99
rect 260 -101 262 -99
rect 286 -101 294 -94
rect 255 -106 262 -101
rect 255 -108 258 -106
rect 260 -108 262 -106
rect 255 -110 262 -108
rect 269 -109 274 -101
rect 255 -122 260 -110
rect 267 -111 274 -109
rect 267 -113 269 -111
rect 271 -113 274 -111
rect 267 -115 274 -113
rect 269 -122 274 -115
rect 276 -122 281 -101
rect 283 -112 294 -101
rect 296 -99 301 -94
rect 296 -101 303 -99
rect 296 -103 299 -101
rect 301 -103 303 -101
rect 336 -102 342 -95
rect 296 -108 303 -103
rect 296 -110 299 -108
rect 301 -110 303 -108
rect 296 -112 303 -110
rect 315 -111 322 -102
rect 283 -118 292 -112
rect 315 -113 317 -111
rect 319 -113 322 -111
rect 315 -115 322 -113
rect 324 -104 332 -102
rect 324 -106 327 -104
rect 329 -106 332 -104
rect 324 -111 332 -106
rect 324 -113 327 -111
rect 329 -113 332 -111
rect 324 -115 332 -113
rect 334 -109 342 -102
rect 334 -111 337 -109
rect 339 -111 342 -109
rect 334 -113 342 -111
rect 344 -97 351 -95
rect 380 -97 385 -94
rect 344 -99 347 -97
rect 349 -99 351 -97
rect 344 -104 351 -99
rect 344 -106 347 -104
rect 349 -106 351 -104
rect 344 -108 351 -106
rect 355 -99 362 -97
rect 355 -101 357 -99
rect 359 -101 362 -99
rect 355 -106 362 -101
rect 355 -108 357 -106
rect 359 -108 362 -106
rect 344 -113 349 -108
rect 355 -110 362 -108
rect 334 -115 340 -113
rect 283 -120 288 -118
rect 290 -120 292 -118
rect 283 -122 292 -120
rect 357 -122 362 -110
rect 364 -110 375 -97
rect 377 -99 385 -97
rect 377 -101 380 -99
rect 382 -101 385 -99
rect 377 -110 385 -101
rect 364 -118 373 -110
rect 364 -120 368 -118
rect 370 -120 373 -118
rect 380 -119 385 -110
rect 387 -119 392 -94
rect 394 -111 410 -94
rect 394 -113 403 -111
rect 405 -113 410 -111
rect 394 -118 410 -113
rect 394 -119 403 -118
rect 364 -122 373 -120
rect 396 -120 403 -119
rect 405 -120 410 -118
rect 396 -122 410 -120
rect 412 -103 420 -94
rect 412 -105 415 -103
rect 417 -105 420 -103
rect 412 -110 420 -105
rect 412 -112 415 -110
rect 417 -112 420 -110
rect 412 -122 420 -112
rect 422 -111 430 -94
rect 422 -113 425 -111
rect 427 -113 430 -111
rect 422 -118 430 -113
rect 422 -120 425 -118
rect 427 -120 430 -118
rect 422 -122 430 -120
rect 432 -96 439 -94
rect 432 -98 435 -96
rect 437 -98 439 -96
rect 432 -103 439 -98
rect 432 -105 435 -103
rect 437 -105 439 -103
rect 432 -107 439 -105
rect 445 -96 452 -94
rect 445 -98 447 -96
rect 449 -98 452 -96
rect 445 -103 452 -98
rect 445 -105 447 -103
rect 449 -105 452 -103
rect 445 -107 452 -105
rect 432 -122 437 -107
rect 447 -122 452 -107
rect 454 -111 462 -94
rect 454 -113 457 -111
rect 459 -113 462 -111
rect 454 -118 462 -113
rect 454 -120 457 -118
rect 459 -120 462 -118
rect 454 -122 462 -120
rect 464 -103 472 -94
rect 464 -105 467 -103
rect 469 -105 472 -103
rect 464 -110 472 -105
rect 464 -112 467 -110
rect 469 -112 472 -110
rect 464 -122 472 -112
rect 474 -111 490 -94
rect 474 -113 479 -111
rect 481 -113 490 -111
rect 474 -118 490 -113
rect 474 -120 479 -118
rect 481 -119 490 -118
rect 492 -119 497 -94
rect 499 -97 504 -94
rect 499 -99 507 -97
rect 499 -101 502 -99
rect 504 -101 507 -99
rect 499 -110 507 -101
rect 509 -110 520 -97
rect 499 -119 504 -110
rect 511 -118 520 -110
rect 481 -120 488 -119
rect 474 -122 488 -120
rect 511 -120 514 -118
rect 516 -120 520 -118
rect 511 -122 520 -120
rect 522 -99 529 -97
rect 522 -101 525 -99
rect 527 -101 529 -99
rect 553 -101 561 -94
rect 522 -106 529 -101
rect 522 -108 525 -106
rect 527 -108 529 -106
rect 522 -110 529 -108
rect 536 -109 541 -101
rect 522 -122 527 -110
rect 534 -111 541 -109
rect 534 -113 536 -111
rect 538 -113 541 -111
rect 534 -115 541 -113
rect 536 -122 541 -115
rect 543 -122 548 -101
rect 550 -112 561 -101
rect 563 -99 568 -94
rect 563 -101 570 -99
rect 563 -103 566 -101
rect 568 -103 570 -101
rect 603 -102 609 -95
rect 563 -108 570 -103
rect 563 -110 566 -108
rect 568 -110 570 -108
rect 563 -112 570 -110
rect 582 -111 589 -102
rect 550 -118 559 -112
rect 582 -113 584 -111
rect 586 -113 589 -111
rect 582 -115 589 -113
rect 591 -104 599 -102
rect 591 -106 594 -104
rect 596 -106 599 -104
rect 591 -111 599 -106
rect 591 -113 594 -111
rect 596 -113 599 -111
rect 591 -115 599 -113
rect 601 -109 609 -102
rect 601 -111 604 -109
rect 606 -111 609 -109
rect 601 -113 609 -111
rect 611 -97 618 -95
rect 647 -97 652 -94
rect 611 -99 614 -97
rect 616 -99 618 -97
rect 611 -104 618 -99
rect 611 -106 614 -104
rect 616 -106 618 -104
rect 611 -108 618 -106
rect 622 -99 629 -97
rect 622 -101 624 -99
rect 626 -101 629 -99
rect 622 -106 629 -101
rect 622 -108 624 -106
rect 626 -108 629 -106
rect 611 -113 616 -108
rect 622 -110 629 -108
rect 601 -115 607 -113
rect 550 -120 555 -118
rect 557 -120 559 -118
rect 550 -122 559 -120
rect 624 -122 629 -110
rect 631 -110 642 -97
rect 644 -99 652 -97
rect 644 -101 647 -99
rect 649 -101 652 -99
rect 644 -110 652 -101
rect 631 -118 640 -110
rect 631 -120 635 -118
rect 637 -120 640 -118
rect 647 -119 652 -110
rect 654 -119 659 -94
rect 661 -111 677 -94
rect 661 -113 670 -111
rect 672 -113 677 -111
rect 661 -118 677 -113
rect 661 -119 670 -118
rect 631 -122 640 -120
rect 663 -120 670 -119
rect 672 -120 677 -118
rect 663 -122 677 -120
rect 679 -103 687 -94
rect 679 -105 682 -103
rect 684 -105 687 -103
rect 679 -110 687 -105
rect 679 -112 682 -110
rect 684 -112 687 -110
rect 679 -122 687 -112
rect 689 -111 697 -94
rect 689 -113 692 -111
rect 694 -113 697 -111
rect 689 -118 697 -113
rect 689 -120 692 -118
rect 694 -120 697 -118
rect 689 -122 697 -120
rect 699 -96 706 -94
rect 699 -98 702 -96
rect 704 -98 706 -96
rect 699 -103 706 -98
rect 699 -105 702 -103
rect 704 -105 706 -103
rect 699 -107 706 -105
rect 712 -96 719 -94
rect 712 -98 714 -96
rect 716 -98 719 -96
rect 712 -103 719 -98
rect 712 -105 714 -103
rect 716 -105 719 -103
rect 712 -107 719 -105
rect 699 -122 704 -107
rect 714 -122 719 -107
rect 721 -111 729 -94
rect 721 -113 724 -111
rect 726 -113 729 -111
rect 721 -118 729 -113
rect 721 -120 724 -118
rect 726 -120 729 -118
rect 721 -122 729 -120
rect 731 -103 739 -94
rect 731 -105 734 -103
rect 736 -105 739 -103
rect 731 -110 739 -105
rect 731 -112 734 -110
rect 736 -112 739 -110
rect 731 -122 739 -112
rect 741 -111 757 -94
rect 741 -113 746 -111
rect 748 -113 757 -111
rect 741 -118 757 -113
rect 741 -120 746 -118
rect 748 -119 757 -118
rect 759 -119 764 -94
rect 766 -97 771 -94
rect 766 -99 774 -97
rect 766 -101 769 -99
rect 771 -101 774 -99
rect 766 -110 774 -101
rect 776 -110 787 -97
rect 766 -119 771 -110
rect 778 -118 787 -110
rect 748 -120 755 -119
rect 741 -122 755 -120
rect 778 -120 781 -118
rect 783 -120 787 -118
rect 778 -122 787 -120
rect 789 -99 796 -97
rect 789 -101 792 -99
rect 794 -101 796 -99
rect 820 -101 828 -94
rect 789 -106 796 -101
rect 789 -108 792 -106
rect 794 -108 796 -106
rect 789 -110 796 -108
rect 803 -109 808 -101
rect 789 -122 794 -110
rect 801 -111 808 -109
rect 801 -113 803 -111
rect 805 -113 808 -111
rect 801 -115 808 -113
rect 803 -122 808 -115
rect 810 -122 815 -101
rect 817 -112 828 -101
rect 830 -99 835 -94
rect 830 -101 837 -99
rect 830 -103 833 -101
rect 835 -103 837 -101
rect 870 -102 876 -95
rect 830 -108 837 -103
rect 830 -110 833 -108
rect 835 -110 837 -108
rect 830 -112 837 -110
rect 849 -111 856 -102
rect 817 -118 826 -112
rect 849 -113 851 -111
rect 853 -113 856 -111
rect 849 -115 856 -113
rect 858 -104 866 -102
rect 858 -106 861 -104
rect 863 -106 866 -104
rect 858 -111 866 -106
rect 858 -113 861 -111
rect 863 -113 866 -111
rect 858 -115 866 -113
rect 868 -109 876 -102
rect 868 -111 871 -109
rect 873 -111 876 -109
rect 868 -113 876 -111
rect 878 -97 885 -95
rect 914 -97 919 -94
rect 878 -99 881 -97
rect 883 -99 885 -97
rect 878 -104 885 -99
rect 878 -106 881 -104
rect 883 -106 885 -104
rect 878 -108 885 -106
rect 889 -99 896 -97
rect 889 -101 891 -99
rect 893 -101 896 -99
rect 889 -106 896 -101
rect 889 -108 891 -106
rect 893 -108 896 -106
rect 878 -113 883 -108
rect 889 -110 896 -108
rect 868 -115 874 -113
rect 817 -120 822 -118
rect 824 -120 826 -118
rect 817 -122 826 -120
rect 891 -122 896 -110
rect 898 -110 909 -97
rect 911 -99 919 -97
rect 911 -101 914 -99
rect 916 -101 919 -99
rect 911 -110 919 -101
rect 898 -118 907 -110
rect 898 -120 902 -118
rect 904 -120 907 -118
rect 914 -119 919 -110
rect 921 -119 926 -94
rect 928 -111 944 -94
rect 928 -113 937 -111
rect 939 -113 944 -111
rect 928 -118 944 -113
rect 928 -119 937 -118
rect 898 -122 907 -120
rect 930 -120 937 -119
rect 939 -120 944 -118
rect 930 -122 944 -120
rect 946 -103 954 -94
rect 946 -105 949 -103
rect 951 -105 954 -103
rect 946 -110 954 -105
rect 946 -112 949 -110
rect 951 -112 954 -110
rect 946 -122 954 -112
rect 956 -111 964 -94
rect 956 -113 959 -111
rect 961 -113 964 -111
rect 956 -118 964 -113
rect 956 -120 959 -118
rect 961 -120 964 -118
rect 956 -122 964 -120
rect 966 -96 973 -94
rect 966 -98 969 -96
rect 971 -98 973 -96
rect 966 -103 973 -98
rect 966 -105 969 -103
rect 971 -105 973 -103
rect 966 -107 973 -105
rect 979 -96 986 -94
rect 979 -98 981 -96
rect 983 -98 986 -96
rect 979 -103 986 -98
rect 979 -105 981 -103
rect 983 -105 986 -103
rect 979 -107 986 -105
rect 966 -122 971 -107
rect 981 -122 986 -107
rect 988 -111 996 -94
rect 988 -113 991 -111
rect 993 -113 996 -111
rect 988 -118 996 -113
rect 988 -120 991 -118
rect 993 -120 996 -118
rect 988 -122 996 -120
rect 998 -103 1006 -94
rect 998 -105 1001 -103
rect 1003 -105 1006 -103
rect 998 -110 1006 -105
rect 998 -112 1001 -110
rect 1003 -112 1006 -110
rect 998 -122 1006 -112
rect 1008 -111 1024 -94
rect 1008 -113 1013 -111
rect 1015 -113 1024 -111
rect 1008 -118 1024 -113
rect 1008 -120 1013 -118
rect 1015 -119 1024 -118
rect 1026 -119 1031 -94
rect 1033 -97 1038 -94
rect 1033 -99 1041 -97
rect 1033 -101 1036 -99
rect 1038 -101 1041 -99
rect 1033 -110 1041 -101
rect 1043 -110 1054 -97
rect 1033 -119 1038 -110
rect 1045 -118 1054 -110
rect 1015 -120 1022 -119
rect 1008 -122 1022 -120
rect 1045 -120 1048 -118
rect 1050 -120 1054 -118
rect 1045 -122 1054 -120
rect 1056 -99 1063 -97
rect 1056 -101 1059 -99
rect 1061 -101 1063 -99
rect 1087 -101 1095 -94
rect 1056 -106 1063 -101
rect 1056 -108 1059 -106
rect 1061 -108 1063 -106
rect 1056 -110 1063 -108
rect 1070 -109 1075 -101
rect 1056 -122 1061 -110
rect 1068 -111 1075 -109
rect 1068 -113 1070 -111
rect 1072 -113 1075 -111
rect 1068 -115 1075 -113
rect 1070 -122 1075 -115
rect 1077 -122 1082 -101
rect 1084 -112 1095 -101
rect 1097 -99 1102 -94
rect 1097 -101 1104 -99
rect 1097 -103 1100 -101
rect 1102 -103 1104 -101
rect 1137 -102 1143 -95
rect 1097 -108 1104 -103
rect 1097 -110 1100 -108
rect 1102 -110 1104 -108
rect 1097 -112 1104 -110
rect 1116 -111 1123 -102
rect 1084 -118 1093 -112
rect 1116 -113 1118 -111
rect 1120 -113 1123 -111
rect 1116 -115 1123 -113
rect 1125 -104 1133 -102
rect 1125 -106 1128 -104
rect 1130 -106 1133 -104
rect 1125 -111 1133 -106
rect 1125 -113 1128 -111
rect 1130 -113 1133 -111
rect 1125 -115 1133 -113
rect 1135 -109 1143 -102
rect 1135 -111 1138 -109
rect 1140 -111 1143 -109
rect 1135 -113 1143 -111
rect 1145 -97 1152 -95
rect 1181 -97 1186 -94
rect 1145 -99 1148 -97
rect 1150 -99 1152 -97
rect 1145 -104 1152 -99
rect 1145 -106 1148 -104
rect 1150 -106 1152 -104
rect 1145 -108 1152 -106
rect 1156 -99 1163 -97
rect 1156 -101 1158 -99
rect 1160 -101 1163 -99
rect 1156 -106 1163 -101
rect 1156 -108 1158 -106
rect 1160 -108 1163 -106
rect 1145 -113 1150 -108
rect 1156 -110 1163 -108
rect 1135 -115 1141 -113
rect 1084 -120 1089 -118
rect 1091 -120 1093 -118
rect 1084 -122 1093 -120
rect 1158 -122 1163 -110
rect 1165 -110 1176 -97
rect 1178 -99 1186 -97
rect 1178 -101 1181 -99
rect 1183 -101 1186 -99
rect 1178 -110 1186 -101
rect 1165 -118 1174 -110
rect 1165 -120 1169 -118
rect 1171 -120 1174 -118
rect 1181 -119 1186 -110
rect 1188 -119 1193 -94
rect 1195 -111 1211 -94
rect 1195 -113 1204 -111
rect 1206 -113 1211 -111
rect 1195 -118 1211 -113
rect 1195 -119 1204 -118
rect 1165 -122 1174 -120
rect 1197 -120 1204 -119
rect 1206 -120 1211 -118
rect 1197 -122 1211 -120
rect 1213 -103 1221 -94
rect 1213 -105 1216 -103
rect 1218 -105 1221 -103
rect 1213 -110 1221 -105
rect 1213 -112 1216 -110
rect 1218 -112 1221 -110
rect 1213 -122 1221 -112
rect 1223 -111 1231 -94
rect 1223 -113 1226 -111
rect 1228 -113 1231 -111
rect 1223 -118 1231 -113
rect 1223 -120 1226 -118
rect 1228 -120 1231 -118
rect 1223 -122 1231 -120
rect 1233 -96 1240 -94
rect 1233 -98 1236 -96
rect 1238 -98 1240 -96
rect 1233 -103 1240 -98
rect 1233 -105 1236 -103
rect 1238 -105 1240 -103
rect 1233 -107 1240 -105
rect 1246 -96 1253 -94
rect 1246 -98 1248 -96
rect 1250 -98 1253 -96
rect 1246 -103 1253 -98
rect 1246 -105 1248 -103
rect 1250 -105 1253 -103
rect 1246 -107 1253 -105
rect 1233 -122 1238 -107
rect 1248 -122 1253 -107
rect 1255 -111 1263 -94
rect 1255 -113 1258 -111
rect 1260 -113 1263 -111
rect 1255 -118 1263 -113
rect 1255 -120 1258 -118
rect 1260 -120 1263 -118
rect 1255 -122 1263 -120
rect 1265 -103 1273 -94
rect 1265 -105 1268 -103
rect 1270 -105 1273 -103
rect 1265 -110 1273 -105
rect 1265 -112 1268 -110
rect 1270 -112 1273 -110
rect 1265 -122 1273 -112
rect 1275 -111 1291 -94
rect 1275 -113 1280 -111
rect 1282 -113 1291 -111
rect 1275 -118 1291 -113
rect 1275 -120 1280 -118
rect 1282 -119 1291 -118
rect 1293 -119 1298 -94
rect 1300 -97 1305 -94
rect 1300 -99 1308 -97
rect 1300 -101 1303 -99
rect 1305 -101 1308 -99
rect 1300 -110 1308 -101
rect 1310 -110 1321 -97
rect 1300 -119 1305 -110
rect 1312 -118 1321 -110
rect 1282 -120 1289 -119
rect 1275 -122 1289 -120
rect 1312 -120 1315 -118
rect 1317 -120 1321 -118
rect 1312 -122 1321 -120
rect 1323 -99 1330 -97
rect 1323 -101 1326 -99
rect 1328 -101 1330 -99
rect 1354 -101 1362 -94
rect 1323 -106 1330 -101
rect 1323 -108 1326 -106
rect 1328 -108 1330 -106
rect 1323 -110 1330 -108
rect 1337 -109 1342 -101
rect 1323 -122 1328 -110
rect 1335 -111 1342 -109
rect 1335 -113 1337 -111
rect 1339 -113 1342 -111
rect 1335 -115 1342 -113
rect 1337 -122 1342 -115
rect 1344 -122 1349 -101
rect 1351 -112 1362 -101
rect 1364 -99 1369 -94
rect 1364 -101 1371 -99
rect 1364 -103 1367 -101
rect 1369 -103 1371 -101
rect 1404 -102 1410 -95
rect 1364 -108 1371 -103
rect 1364 -110 1367 -108
rect 1369 -110 1371 -108
rect 1364 -112 1371 -110
rect 1383 -111 1390 -102
rect 1351 -118 1360 -112
rect 1383 -113 1385 -111
rect 1387 -113 1390 -111
rect 1383 -115 1390 -113
rect 1392 -104 1400 -102
rect 1392 -106 1395 -104
rect 1397 -106 1400 -104
rect 1392 -111 1400 -106
rect 1392 -113 1395 -111
rect 1397 -113 1400 -111
rect 1392 -115 1400 -113
rect 1402 -109 1410 -102
rect 1402 -111 1405 -109
rect 1407 -111 1410 -109
rect 1402 -113 1410 -111
rect 1412 -97 1419 -95
rect 1448 -97 1453 -94
rect 1412 -99 1415 -97
rect 1417 -99 1419 -97
rect 1412 -104 1419 -99
rect 1412 -106 1415 -104
rect 1417 -106 1419 -104
rect 1412 -108 1419 -106
rect 1423 -99 1430 -97
rect 1423 -101 1425 -99
rect 1427 -101 1430 -99
rect 1423 -106 1430 -101
rect 1423 -108 1425 -106
rect 1427 -108 1430 -106
rect 1412 -113 1417 -108
rect 1423 -110 1430 -108
rect 1402 -115 1408 -113
rect 1351 -120 1356 -118
rect 1358 -120 1360 -118
rect 1351 -122 1360 -120
rect 1425 -122 1430 -110
rect 1432 -110 1443 -97
rect 1445 -99 1453 -97
rect 1445 -101 1448 -99
rect 1450 -101 1453 -99
rect 1445 -110 1453 -101
rect 1432 -118 1441 -110
rect 1432 -120 1436 -118
rect 1438 -120 1441 -118
rect 1448 -119 1453 -110
rect 1455 -119 1460 -94
rect 1462 -111 1478 -94
rect 1462 -113 1471 -111
rect 1473 -113 1478 -111
rect 1462 -118 1478 -113
rect 1462 -119 1471 -118
rect 1432 -122 1441 -120
rect 1464 -120 1471 -119
rect 1473 -120 1478 -118
rect 1464 -122 1478 -120
rect 1480 -103 1488 -94
rect 1480 -105 1483 -103
rect 1485 -105 1488 -103
rect 1480 -110 1488 -105
rect 1480 -112 1483 -110
rect 1485 -112 1488 -110
rect 1480 -122 1488 -112
rect 1490 -111 1498 -94
rect 1490 -113 1493 -111
rect 1495 -113 1498 -111
rect 1490 -118 1498 -113
rect 1490 -120 1493 -118
rect 1495 -120 1498 -118
rect 1490 -122 1498 -120
rect 1500 -96 1507 -94
rect 1500 -98 1503 -96
rect 1505 -98 1507 -96
rect 1500 -103 1507 -98
rect 1500 -105 1503 -103
rect 1505 -105 1507 -103
rect 1500 -107 1507 -105
rect 1513 -96 1520 -94
rect 1513 -98 1515 -96
rect 1517 -98 1520 -96
rect 1513 -103 1520 -98
rect 1513 -105 1515 -103
rect 1517 -105 1520 -103
rect 1513 -107 1520 -105
rect 1500 -122 1505 -107
rect 1515 -122 1520 -107
rect 1522 -111 1530 -94
rect 1522 -113 1525 -111
rect 1527 -113 1530 -111
rect 1522 -118 1530 -113
rect 1522 -120 1525 -118
rect 1527 -120 1530 -118
rect 1522 -122 1530 -120
rect 1532 -103 1540 -94
rect 1532 -105 1535 -103
rect 1537 -105 1540 -103
rect 1532 -110 1540 -105
rect 1532 -112 1535 -110
rect 1537 -112 1540 -110
rect 1532 -122 1540 -112
rect 1542 -111 1558 -94
rect 1542 -113 1547 -111
rect 1549 -113 1558 -111
rect 1542 -118 1558 -113
rect 1542 -120 1547 -118
rect 1549 -119 1558 -118
rect 1560 -119 1565 -94
rect 1567 -97 1572 -94
rect 1567 -99 1575 -97
rect 1567 -101 1570 -99
rect 1572 -101 1575 -99
rect 1567 -110 1575 -101
rect 1577 -110 1588 -97
rect 1567 -119 1572 -110
rect 1579 -118 1588 -110
rect 1549 -120 1556 -119
rect 1542 -122 1556 -120
rect 1579 -120 1582 -118
rect 1584 -120 1588 -118
rect 1579 -122 1588 -120
rect 1590 -99 1597 -97
rect 1590 -101 1593 -99
rect 1595 -101 1597 -99
rect 1621 -101 1629 -94
rect 1590 -106 1597 -101
rect 1590 -108 1593 -106
rect 1595 -108 1597 -106
rect 1590 -110 1597 -108
rect 1604 -109 1609 -101
rect 1590 -122 1595 -110
rect 1602 -111 1609 -109
rect 1602 -113 1604 -111
rect 1606 -113 1609 -111
rect 1602 -115 1609 -113
rect 1604 -122 1609 -115
rect 1611 -122 1616 -101
rect 1618 -112 1629 -101
rect 1631 -99 1636 -94
rect 1631 -101 1638 -99
rect 1631 -103 1634 -101
rect 1636 -103 1638 -101
rect 1671 -102 1677 -95
rect 1631 -108 1638 -103
rect 1631 -110 1634 -108
rect 1636 -110 1638 -108
rect 1631 -112 1638 -110
rect 1650 -111 1657 -102
rect 1618 -118 1627 -112
rect 1650 -113 1652 -111
rect 1654 -113 1657 -111
rect 1650 -115 1657 -113
rect 1659 -104 1667 -102
rect 1659 -106 1662 -104
rect 1664 -106 1667 -104
rect 1659 -111 1667 -106
rect 1659 -113 1662 -111
rect 1664 -113 1667 -111
rect 1659 -115 1667 -113
rect 1669 -109 1677 -102
rect 1669 -111 1672 -109
rect 1674 -111 1677 -109
rect 1669 -113 1677 -111
rect 1679 -97 1686 -95
rect 1715 -97 1720 -94
rect 1679 -99 1682 -97
rect 1684 -99 1686 -97
rect 1679 -104 1686 -99
rect 1679 -106 1682 -104
rect 1684 -106 1686 -104
rect 1679 -108 1686 -106
rect 1690 -99 1697 -97
rect 1690 -101 1692 -99
rect 1694 -101 1697 -99
rect 1690 -106 1697 -101
rect 1690 -108 1692 -106
rect 1694 -108 1697 -106
rect 1679 -113 1684 -108
rect 1690 -110 1697 -108
rect 1669 -115 1675 -113
rect 1618 -120 1623 -118
rect 1625 -120 1627 -118
rect 1618 -122 1627 -120
rect 1692 -122 1697 -110
rect 1699 -110 1710 -97
rect 1712 -99 1720 -97
rect 1712 -101 1715 -99
rect 1717 -101 1720 -99
rect 1712 -110 1720 -101
rect 1699 -118 1708 -110
rect 1699 -120 1703 -118
rect 1705 -120 1708 -118
rect 1715 -119 1720 -110
rect 1722 -119 1727 -94
rect 1729 -111 1745 -94
rect 1729 -113 1738 -111
rect 1740 -113 1745 -111
rect 1729 -118 1745 -113
rect 1729 -119 1738 -118
rect 1699 -122 1708 -120
rect 1731 -120 1738 -119
rect 1740 -120 1745 -118
rect 1731 -122 1745 -120
rect 1747 -103 1755 -94
rect 1747 -105 1750 -103
rect 1752 -105 1755 -103
rect 1747 -110 1755 -105
rect 1747 -112 1750 -110
rect 1752 -112 1755 -110
rect 1747 -122 1755 -112
rect 1757 -111 1765 -94
rect 1757 -113 1760 -111
rect 1762 -113 1765 -111
rect 1757 -118 1765 -113
rect 1757 -120 1760 -118
rect 1762 -120 1765 -118
rect 1757 -122 1765 -120
rect 1767 -96 1774 -94
rect 1767 -98 1770 -96
rect 1772 -98 1774 -96
rect 1767 -103 1774 -98
rect 1767 -105 1770 -103
rect 1772 -105 1774 -103
rect 1767 -107 1774 -105
rect 1780 -96 1787 -94
rect 1780 -98 1782 -96
rect 1784 -98 1787 -96
rect 1780 -103 1787 -98
rect 1780 -105 1782 -103
rect 1784 -105 1787 -103
rect 1780 -107 1787 -105
rect 1767 -122 1772 -107
rect 1782 -122 1787 -107
rect 1789 -111 1797 -94
rect 1789 -113 1792 -111
rect 1794 -113 1797 -111
rect 1789 -118 1797 -113
rect 1789 -120 1792 -118
rect 1794 -120 1797 -118
rect 1789 -122 1797 -120
rect 1799 -103 1807 -94
rect 1799 -105 1802 -103
rect 1804 -105 1807 -103
rect 1799 -110 1807 -105
rect 1799 -112 1802 -110
rect 1804 -112 1807 -110
rect 1799 -122 1807 -112
rect 1809 -111 1825 -94
rect 1809 -113 1814 -111
rect 1816 -113 1825 -111
rect 1809 -118 1825 -113
rect 1809 -120 1814 -118
rect 1816 -119 1825 -118
rect 1827 -119 1832 -94
rect 1834 -97 1839 -94
rect 1834 -99 1842 -97
rect 1834 -101 1837 -99
rect 1839 -101 1842 -99
rect 1834 -110 1842 -101
rect 1844 -110 1855 -97
rect 1834 -119 1839 -110
rect 1846 -118 1855 -110
rect 1816 -120 1823 -119
rect 1809 -122 1823 -120
rect 1846 -120 1849 -118
rect 1851 -120 1855 -118
rect 1846 -122 1855 -120
rect 1857 -99 1864 -97
rect 1857 -101 1860 -99
rect 1862 -101 1864 -99
rect 1888 -101 1896 -94
rect 1857 -106 1864 -101
rect 1857 -108 1860 -106
rect 1862 -108 1864 -106
rect 1857 -110 1864 -108
rect 1871 -109 1876 -101
rect 1857 -122 1862 -110
rect 1869 -111 1876 -109
rect 1869 -113 1871 -111
rect 1873 -113 1876 -111
rect 1869 -115 1876 -113
rect 1871 -122 1876 -115
rect 1878 -122 1883 -101
rect 1885 -112 1896 -101
rect 1898 -99 1903 -94
rect 1920 -97 1927 -95
rect 1920 -99 1922 -97
rect 1924 -99 1927 -97
rect 1898 -101 1905 -99
rect 1920 -101 1927 -99
rect 1898 -103 1901 -101
rect 1903 -103 1905 -101
rect 1898 -108 1905 -103
rect 1898 -110 1901 -108
rect 1903 -110 1905 -108
rect 1898 -112 1905 -110
rect 1885 -118 1894 -112
rect 1885 -120 1890 -118
rect 1892 -120 1894 -118
rect 1885 -122 1894 -120
rect 1922 -122 1927 -101
rect 1929 -111 1943 -95
rect 1929 -113 1932 -111
rect 1934 -113 1943 -111
rect 1945 -97 1953 -95
rect 1945 -99 1948 -97
rect 1950 -99 1953 -97
rect 1945 -104 1953 -99
rect 1945 -106 1948 -104
rect 1950 -106 1953 -104
rect 1945 -113 1953 -106
rect 1955 -104 1963 -95
rect 1955 -106 1958 -104
rect 1960 -106 1963 -104
rect 1955 -113 1963 -106
rect 1929 -118 1941 -113
rect 1929 -120 1932 -118
rect 1934 -120 1941 -118
rect 1929 -122 1941 -120
rect 1958 -122 1963 -113
rect 1965 -110 1970 -95
rect 2001 -97 2006 -94
rect 1976 -99 1983 -97
rect 1976 -101 1978 -99
rect 1980 -101 1983 -99
rect 1976 -106 1983 -101
rect 1976 -108 1978 -106
rect 1980 -108 1983 -106
rect 1976 -110 1983 -108
rect 1965 -112 1972 -110
rect 1965 -114 1968 -112
rect 1970 -114 1972 -112
rect 1965 -116 1972 -114
rect 1965 -122 1970 -116
rect 1978 -122 1983 -110
rect 1985 -110 1996 -97
rect 1998 -99 2006 -97
rect 1998 -101 2001 -99
rect 2003 -101 2006 -99
rect 1998 -110 2006 -101
rect 1985 -118 1994 -110
rect 1985 -120 1989 -118
rect 1991 -120 1994 -118
rect 2001 -119 2006 -110
rect 2008 -119 2013 -94
rect 2015 -111 2031 -94
rect 2015 -113 2024 -111
rect 2026 -113 2031 -111
rect 2015 -118 2031 -113
rect 2015 -119 2024 -118
rect 1985 -122 1994 -120
rect 2017 -120 2024 -119
rect 2026 -120 2031 -118
rect 2017 -122 2031 -120
rect 2033 -103 2041 -94
rect 2033 -105 2036 -103
rect 2038 -105 2041 -103
rect 2033 -110 2041 -105
rect 2033 -112 2036 -110
rect 2038 -112 2041 -110
rect 2033 -122 2041 -112
rect 2043 -111 2051 -94
rect 2043 -113 2046 -111
rect 2048 -113 2051 -111
rect 2043 -118 2051 -113
rect 2043 -120 2046 -118
rect 2048 -120 2051 -118
rect 2043 -122 2051 -120
rect 2053 -96 2060 -94
rect 2053 -98 2056 -96
rect 2058 -98 2060 -96
rect 2053 -103 2060 -98
rect 2053 -105 2056 -103
rect 2058 -105 2060 -103
rect 2053 -107 2060 -105
rect 2066 -96 2073 -94
rect 2066 -98 2068 -96
rect 2070 -98 2073 -96
rect 2066 -103 2073 -98
rect 2066 -105 2068 -103
rect 2070 -105 2073 -103
rect 2066 -107 2073 -105
rect 2053 -122 2058 -107
rect 2068 -122 2073 -107
rect 2075 -111 2083 -94
rect 2075 -113 2078 -111
rect 2080 -113 2083 -111
rect 2075 -118 2083 -113
rect 2075 -120 2078 -118
rect 2080 -120 2083 -118
rect 2075 -122 2083 -120
rect 2085 -103 2093 -94
rect 2085 -105 2088 -103
rect 2090 -105 2093 -103
rect 2085 -110 2093 -105
rect 2085 -112 2088 -110
rect 2090 -112 2093 -110
rect 2085 -122 2093 -112
rect 2095 -111 2111 -94
rect 2095 -113 2100 -111
rect 2102 -113 2111 -111
rect 2095 -118 2111 -113
rect 2095 -120 2100 -118
rect 2102 -119 2111 -118
rect 2113 -119 2118 -94
rect 2120 -97 2125 -94
rect 2120 -99 2128 -97
rect 2120 -101 2123 -99
rect 2125 -101 2128 -99
rect 2120 -110 2128 -101
rect 2130 -110 2141 -97
rect 2120 -119 2125 -110
rect 2132 -118 2141 -110
rect 2102 -120 2109 -119
rect 2095 -122 2109 -120
rect 2132 -120 2135 -118
rect 2137 -120 2141 -118
rect 2132 -122 2141 -120
rect 2143 -99 2150 -97
rect 2143 -101 2146 -99
rect 2148 -101 2150 -99
rect 2174 -101 2182 -94
rect 2143 -106 2150 -101
rect 2143 -108 2146 -106
rect 2148 -108 2150 -106
rect 2143 -110 2150 -108
rect 2157 -109 2162 -101
rect 2143 -122 2148 -110
rect 2155 -111 2162 -109
rect 2155 -113 2157 -111
rect 2159 -113 2162 -111
rect 2155 -115 2162 -113
rect 2157 -122 2162 -115
rect 2164 -122 2169 -101
rect 2171 -112 2182 -101
rect 2184 -99 2189 -94
rect 2199 -96 2206 -94
rect 2199 -98 2201 -96
rect 2203 -98 2206 -96
rect 2184 -101 2191 -99
rect 2199 -100 2206 -98
rect 2184 -103 2187 -101
rect 2189 -103 2191 -101
rect 2201 -102 2206 -100
rect 2208 -102 2214 -94
rect 2184 -108 2191 -103
rect 2184 -110 2187 -108
rect 2189 -110 2191 -108
rect 2184 -112 2191 -110
rect 2210 -106 2214 -102
rect 2267 -96 2274 -94
rect 2267 -98 2269 -96
rect 2271 -98 2274 -96
rect 2267 -100 2274 -98
rect 2269 -102 2274 -100
rect 2276 -102 2282 -94
rect 2245 -106 2250 -104
rect 2210 -110 2216 -106
rect 2171 -118 2180 -112
rect 2171 -120 2176 -118
rect 2178 -120 2180 -118
rect 2209 -118 2216 -110
rect 2171 -122 2180 -120
rect 2209 -120 2211 -118
rect 2213 -120 2216 -118
rect 2209 -122 2216 -120
rect 2218 -122 2223 -106
rect 2225 -108 2233 -106
rect 2225 -110 2228 -108
rect 2230 -110 2233 -108
rect 2225 -122 2233 -110
rect 2235 -122 2240 -106
rect 2242 -118 2250 -106
rect 2242 -120 2245 -118
rect 2247 -120 2250 -118
rect 2242 -122 2250 -120
rect 2252 -109 2257 -104
rect 2278 -106 2282 -102
rect 2313 -106 2318 -104
rect 2252 -111 2259 -109
rect 2278 -110 2284 -106
rect 2252 -113 2255 -111
rect 2257 -113 2259 -111
rect 2252 -115 2259 -113
rect 2252 -122 2257 -115
rect 2277 -118 2284 -110
rect 2277 -120 2279 -118
rect 2281 -120 2284 -118
rect 2277 -122 2284 -120
rect 2286 -122 2291 -106
rect 2293 -108 2301 -106
rect 2293 -110 2296 -108
rect 2298 -110 2301 -108
rect 2293 -122 2301 -110
rect 2303 -122 2308 -106
rect 2310 -118 2318 -106
rect 2310 -120 2313 -118
rect 2315 -120 2318 -118
rect 2310 -122 2318 -120
rect 2320 -109 2325 -104
rect 2320 -111 2327 -109
rect 2320 -113 2323 -111
rect 2325 -113 2327 -111
rect 2320 -115 2327 -113
rect 2320 -122 2325 -115
rect 8 -143 15 -141
rect 8 -145 10 -143
rect 12 -145 15 -143
rect 8 -154 15 -145
rect 17 -143 25 -141
rect 17 -145 20 -143
rect 22 -145 25 -143
rect 17 -150 25 -145
rect 17 -152 20 -150
rect 22 -152 25 -150
rect 17 -154 25 -152
rect 27 -143 33 -141
rect 48 -143 55 -141
rect 27 -145 35 -143
rect 27 -147 30 -145
rect 32 -147 35 -145
rect 27 -154 35 -147
rect 29 -161 35 -154
rect 37 -145 42 -143
rect 48 -145 50 -143
rect 52 -145 55 -143
rect 37 -147 44 -145
rect 37 -149 40 -147
rect 42 -149 44 -147
rect 37 -155 44 -149
rect 48 -154 55 -145
rect 57 -143 65 -141
rect 57 -145 60 -143
rect 62 -145 65 -143
rect 57 -150 65 -145
rect 57 -152 60 -150
rect 62 -152 65 -150
rect 57 -154 65 -152
rect 67 -143 73 -141
rect 67 -145 75 -143
rect 67 -147 70 -145
rect 72 -147 75 -145
rect 67 -154 75 -147
rect 37 -157 40 -155
rect 42 -157 44 -155
rect 37 -161 44 -157
rect 69 -161 75 -154
rect 77 -148 82 -143
rect 90 -146 95 -134
rect 88 -148 95 -146
rect 77 -150 84 -148
rect 77 -152 80 -150
rect 82 -152 84 -150
rect 77 -157 84 -152
rect 77 -159 80 -157
rect 82 -159 84 -157
rect 88 -150 90 -148
rect 92 -150 95 -148
rect 88 -155 95 -150
rect 88 -157 90 -155
rect 92 -157 95 -155
rect 88 -159 95 -157
rect 97 -136 106 -134
rect 97 -138 101 -136
rect 103 -138 106 -136
rect 129 -136 143 -134
rect 129 -137 136 -136
rect 97 -146 106 -138
rect 113 -146 118 -137
rect 97 -159 108 -146
rect 110 -155 118 -146
rect 110 -157 113 -155
rect 115 -157 118 -155
rect 110 -159 118 -157
rect 77 -161 84 -159
rect 113 -162 118 -159
rect 120 -162 125 -137
rect 127 -138 136 -137
rect 138 -138 143 -136
rect 127 -143 143 -138
rect 127 -145 136 -143
rect 138 -145 143 -143
rect 127 -162 143 -145
rect 145 -144 153 -134
rect 145 -146 148 -144
rect 150 -146 153 -144
rect 145 -151 153 -146
rect 145 -153 148 -151
rect 150 -153 153 -151
rect 145 -162 153 -153
rect 155 -136 163 -134
rect 155 -138 158 -136
rect 160 -138 163 -136
rect 155 -143 163 -138
rect 155 -145 158 -143
rect 160 -145 163 -143
rect 155 -162 163 -145
rect 165 -149 170 -134
rect 180 -149 185 -134
rect 165 -151 172 -149
rect 165 -153 168 -151
rect 170 -153 172 -151
rect 165 -158 172 -153
rect 165 -160 168 -158
rect 170 -160 172 -158
rect 165 -162 172 -160
rect 178 -151 185 -149
rect 178 -153 180 -151
rect 182 -153 185 -151
rect 178 -158 185 -153
rect 178 -160 180 -158
rect 182 -160 185 -158
rect 178 -162 185 -160
rect 187 -136 195 -134
rect 187 -138 190 -136
rect 192 -138 195 -136
rect 187 -143 195 -138
rect 187 -145 190 -143
rect 192 -145 195 -143
rect 187 -162 195 -145
rect 197 -144 205 -134
rect 197 -146 200 -144
rect 202 -146 205 -144
rect 197 -151 205 -146
rect 197 -153 200 -151
rect 202 -153 205 -151
rect 197 -162 205 -153
rect 207 -136 221 -134
rect 207 -138 212 -136
rect 214 -137 221 -136
rect 244 -136 253 -134
rect 214 -138 223 -137
rect 207 -143 223 -138
rect 207 -145 212 -143
rect 214 -145 223 -143
rect 207 -162 223 -145
rect 225 -162 230 -137
rect 232 -146 237 -137
rect 244 -138 247 -136
rect 249 -138 253 -136
rect 244 -146 253 -138
rect 232 -155 240 -146
rect 232 -157 235 -155
rect 237 -157 240 -155
rect 232 -159 240 -157
rect 242 -159 253 -146
rect 255 -146 260 -134
rect 269 -141 274 -134
rect 267 -143 274 -141
rect 267 -145 269 -143
rect 271 -145 274 -143
rect 255 -148 262 -146
rect 267 -147 274 -145
rect 255 -150 258 -148
rect 260 -150 262 -148
rect 255 -155 262 -150
rect 269 -155 274 -147
rect 276 -155 281 -134
rect 283 -136 292 -134
rect 283 -138 288 -136
rect 290 -138 292 -136
rect 283 -144 292 -138
rect 315 -143 322 -141
rect 283 -155 294 -144
rect 255 -157 258 -155
rect 260 -157 262 -155
rect 255 -159 262 -157
rect 232 -162 237 -159
rect 286 -162 294 -155
rect 296 -146 303 -144
rect 296 -148 299 -146
rect 301 -148 303 -146
rect 296 -153 303 -148
rect 296 -155 299 -153
rect 301 -155 303 -153
rect 315 -145 317 -143
rect 319 -145 322 -143
rect 315 -154 322 -145
rect 324 -143 332 -141
rect 324 -145 327 -143
rect 329 -145 332 -143
rect 324 -150 332 -145
rect 324 -152 327 -150
rect 329 -152 332 -150
rect 324 -154 332 -152
rect 334 -143 340 -141
rect 334 -145 342 -143
rect 334 -147 337 -145
rect 339 -147 342 -145
rect 334 -154 342 -147
rect 296 -157 303 -155
rect 296 -162 301 -157
rect 336 -161 342 -154
rect 344 -148 349 -143
rect 357 -146 362 -134
rect 355 -148 362 -146
rect 344 -150 351 -148
rect 344 -152 347 -150
rect 349 -152 351 -150
rect 344 -157 351 -152
rect 344 -159 347 -157
rect 349 -159 351 -157
rect 355 -150 357 -148
rect 359 -150 362 -148
rect 355 -155 362 -150
rect 355 -157 357 -155
rect 359 -157 362 -155
rect 355 -159 362 -157
rect 364 -136 373 -134
rect 364 -138 368 -136
rect 370 -138 373 -136
rect 396 -136 410 -134
rect 396 -137 403 -136
rect 364 -146 373 -138
rect 380 -146 385 -137
rect 364 -159 375 -146
rect 377 -155 385 -146
rect 377 -157 380 -155
rect 382 -157 385 -155
rect 377 -159 385 -157
rect 344 -161 351 -159
rect 380 -162 385 -159
rect 387 -162 392 -137
rect 394 -138 403 -137
rect 405 -138 410 -136
rect 394 -143 410 -138
rect 394 -145 403 -143
rect 405 -145 410 -143
rect 394 -162 410 -145
rect 412 -144 420 -134
rect 412 -146 415 -144
rect 417 -146 420 -144
rect 412 -151 420 -146
rect 412 -153 415 -151
rect 417 -153 420 -151
rect 412 -162 420 -153
rect 422 -136 430 -134
rect 422 -138 425 -136
rect 427 -138 430 -136
rect 422 -143 430 -138
rect 422 -145 425 -143
rect 427 -145 430 -143
rect 422 -162 430 -145
rect 432 -149 437 -134
rect 447 -149 452 -134
rect 432 -151 439 -149
rect 432 -153 435 -151
rect 437 -153 439 -151
rect 432 -158 439 -153
rect 432 -160 435 -158
rect 437 -160 439 -158
rect 432 -162 439 -160
rect 445 -151 452 -149
rect 445 -153 447 -151
rect 449 -153 452 -151
rect 445 -158 452 -153
rect 445 -160 447 -158
rect 449 -160 452 -158
rect 445 -162 452 -160
rect 454 -136 462 -134
rect 454 -138 457 -136
rect 459 -138 462 -136
rect 454 -143 462 -138
rect 454 -145 457 -143
rect 459 -145 462 -143
rect 454 -162 462 -145
rect 464 -144 472 -134
rect 464 -146 467 -144
rect 469 -146 472 -144
rect 464 -151 472 -146
rect 464 -153 467 -151
rect 469 -153 472 -151
rect 464 -162 472 -153
rect 474 -136 488 -134
rect 474 -138 479 -136
rect 481 -137 488 -136
rect 511 -136 520 -134
rect 481 -138 490 -137
rect 474 -143 490 -138
rect 474 -145 479 -143
rect 481 -145 490 -143
rect 474 -162 490 -145
rect 492 -162 497 -137
rect 499 -146 504 -137
rect 511 -138 514 -136
rect 516 -138 520 -136
rect 511 -146 520 -138
rect 499 -155 507 -146
rect 499 -157 502 -155
rect 504 -157 507 -155
rect 499 -159 507 -157
rect 509 -159 520 -146
rect 522 -146 527 -134
rect 536 -141 541 -134
rect 534 -143 541 -141
rect 534 -145 536 -143
rect 538 -145 541 -143
rect 522 -148 529 -146
rect 534 -147 541 -145
rect 522 -150 525 -148
rect 527 -150 529 -148
rect 522 -155 529 -150
rect 536 -155 541 -147
rect 543 -155 548 -134
rect 550 -136 559 -134
rect 550 -138 555 -136
rect 557 -138 559 -136
rect 550 -144 559 -138
rect 582 -143 589 -141
rect 550 -155 561 -144
rect 522 -157 525 -155
rect 527 -157 529 -155
rect 522 -159 529 -157
rect 499 -162 504 -159
rect 553 -162 561 -155
rect 563 -146 570 -144
rect 563 -148 566 -146
rect 568 -148 570 -146
rect 563 -153 570 -148
rect 563 -155 566 -153
rect 568 -155 570 -153
rect 582 -145 584 -143
rect 586 -145 589 -143
rect 582 -154 589 -145
rect 591 -143 599 -141
rect 591 -145 594 -143
rect 596 -145 599 -143
rect 591 -150 599 -145
rect 591 -152 594 -150
rect 596 -152 599 -150
rect 591 -154 599 -152
rect 601 -143 607 -141
rect 601 -145 609 -143
rect 601 -147 604 -145
rect 606 -147 609 -145
rect 601 -154 609 -147
rect 563 -157 570 -155
rect 563 -162 568 -157
rect 603 -161 609 -154
rect 611 -148 616 -143
rect 624 -146 629 -134
rect 622 -148 629 -146
rect 611 -150 618 -148
rect 611 -152 614 -150
rect 616 -152 618 -150
rect 611 -157 618 -152
rect 611 -159 614 -157
rect 616 -159 618 -157
rect 622 -150 624 -148
rect 626 -150 629 -148
rect 622 -155 629 -150
rect 622 -157 624 -155
rect 626 -157 629 -155
rect 622 -159 629 -157
rect 631 -136 640 -134
rect 631 -138 635 -136
rect 637 -138 640 -136
rect 663 -136 677 -134
rect 663 -137 670 -136
rect 631 -146 640 -138
rect 647 -146 652 -137
rect 631 -159 642 -146
rect 644 -155 652 -146
rect 644 -157 647 -155
rect 649 -157 652 -155
rect 644 -159 652 -157
rect 611 -161 618 -159
rect 647 -162 652 -159
rect 654 -162 659 -137
rect 661 -138 670 -137
rect 672 -138 677 -136
rect 661 -143 677 -138
rect 661 -145 670 -143
rect 672 -145 677 -143
rect 661 -162 677 -145
rect 679 -144 687 -134
rect 679 -146 682 -144
rect 684 -146 687 -144
rect 679 -151 687 -146
rect 679 -153 682 -151
rect 684 -153 687 -151
rect 679 -162 687 -153
rect 689 -136 697 -134
rect 689 -138 692 -136
rect 694 -138 697 -136
rect 689 -143 697 -138
rect 689 -145 692 -143
rect 694 -145 697 -143
rect 689 -162 697 -145
rect 699 -149 704 -134
rect 714 -149 719 -134
rect 699 -151 706 -149
rect 699 -153 702 -151
rect 704 -153 706 -151
rect 699 -158 706 -153
rect 699 -160 702 -158
rect 704 -160 706 -158
rect 699 -162 706 -160
rect 712 -151 719 -149
rect 712 -153 714 -151
rect 716 -153 719 -151
rect 712 -158 719 -153
rect 712 -160 714 -158
rect 716 -160 719 -158
rect 712 -162 719 -160
rect 721 -136 729 -134
rect 721 -138 724 -136
rect 726 -138 729 -136
rect 721 -143 729 -138
rect 721 -145 724 -143
rect 726 -145 729 -143
rect 721 -162 729 -145
rect 731 -144 739 -134
rect 731 -146 734 -144
rect 736 -146 739 -144
rect 731 -151 739 -146
rect 731 -153 734 -151
rect 736 -153 739 -151
rect 731 -162 739 -153
rect 741 -136 755 -134
rect 741 -138 746 -136
rect 748 -137 755 -136
rect 778 -136 787 -134
rect 748 -138 757 -137
rect 741 -143 757 -138
rect 741 -145 746 -143
rect 748 -145 757 -143
rect 741 -162 757 -145
rect 759 -162 764 -137
rect 766 -146 771 -137
rect 778 -138 781 -136
rect 783 -138 787 -136
rect 778 -146 787 -138
rect 766 -155 774 -146
rect 766 -157 769 -155
rect 771 -157 774 -155
rect 766 -159 774 -157
rect 776 -159 787 -146
rect 789 -146 794 -134
rect 803 -141 808 -134
rect 801 -143 808 -141
rect 801 -145 803 -143
rect 805 -145 808 -143
rect 789 -148 796 -146
rect 801 -147 808 -145
rect 789 -150 792 -148
rect 794 -150 796 -148
rect 789 -155 796 -150
rect 803 -155 808 -147
rect 810 -155 815 -134
rect 817 -136 826 -134
rect 817 -138 822 -136
rect 824 -138 826 -136
rect 817 -144 826 -138
rect 849 -143 856 -141
rect 817 -155 828 -144
rect 789 -157 792 -155
rect 794 -157 796 -155
rect 789 -159 796 -157
rect 766 -162 771 -159
rect 820 -162 828 -155
rect 830 -146 837 -144
rect 830 -148 833 -146
rect 835 -148 837 -146
rect 830 -153 837 -148
rect 830 -155 833 -153
rect 835 -155 837 -153
rect 849 -145 851 -143
rect 853 -145 856 -143
rect 849 -154 856 -145
rect 858 -143 866 -141
rect 858 -145 861 -143
rect 863 -145 866 -143
rect 858 -150 866 -145
rect 858 -152 861 -150
rect 863 -152 866 -150
rect 858 -154 866 -152
rect 868 -143 874 -141
rect 868 -145 876 -143
rect 868 -147 871 -145
rect 873 -147 876 -145
rect 868 -154 876 -147
rect 830 -157 837 -155
rect 830 -162 835 -157
rect 870 -161 876 -154
rect 878 -148 883 -143
rect 891 -146 896 -134
rect 889 -148 896 -146
rect 878 -150 885 -148
rect 878 -152 881 -150
rect 883 -152 885 -150
rect 878 -157 885 -152
rect 878 -159 881 -157
rect 883 -159 885 -157
rect 889 -150 891 -148
rect 893 -150 896 -148
rect 889 -155 896 -150
rect 889 -157 891 -155
rect 893 -157 896 -155
rect 889 -159 896 -157
rect 898 -136 907 -134
rect 898 -138 902 -136
rect 904 -138 907 -136
rect 930 -136 944 -134
rect 930 -137 937 -136
rect 898 -146 907 -138
rect 914 -146 919 -137
rect 898 -159 909 -146
rect 911 -155 919 -146
rect 911 -157 914 -155
rect 916 -157 919 -155
rect 911 -159 919 -157
rect 878 -161 885 -159
rect 914 -162 919 -159
rect 921 -162 926 -137
rect 928 -138 937 -137
rect 939 -138 944 -136
rect 928 -143 944 -138
rect 928 -145 937 -143
rect 939 -145 944 -143
rect 928 -162 944 -145
rect 946 -144 954 -134
rect 946 -146 949 -144
rect 951 -146 954 -144
rect 946 -151 954 -146
rect 946 -153 949 -151
rect 951 -153 954 -151
rect 946 -162 954 -153
rect 956 -136 964 -134
rect 956 -138 959 -136
rect 961 -138 964 -136
rect 956 -143 964 -138
rect 956 -145 959 -143
rect 961 -145 964 -143
rect 956 -162 964 -145
rect 966 -149 971 -134
rect 981 -149 986 -134
rect 966 -151 973 -149
rect 966 -153 969 -151
rect 971 -153 973 -151
rect 966 -158 973 -153
rect 966 -160 969 -158
rect 971 -160 973 -158
rect 966 -162 973 -160
rect 979 -151 986 -149
rect 979 -153 981 -151
rect 983 -153 986 -151
rect 979 -158 986 -153
rect 979 -160 981 -158
rect 983 -160 986 -158
rect 979 -162 986 -160
rect 988 -136 996 -134
rect 988 -138 991 -136
rect 993 -138 996 -136
rect 988 -143 996 -138
rect 988 -145 991 -143
rect 993 -145 996 -143
rect 988 -162 996 -145
rect 998 -144 1006 -134
rect 998 -146 1001 -144
rect 1003 -146 1006 -144
rect 998 -151 1006 -146
rect 998 -153 1001 -151
rect 1003 -153 1006 -151
rect 998 -162 1006 -153
rect 1008 -136 1022 -134
rect 1008 -138 1013 -136
rect 1015 -137 1022 -136
rect 1045 -136 1054 -134
rect 1015 -138 1024 -137
rect 1008 -143 1024 -138
rect 1008 -145 1013 -143
rect 1015 -145 1024 -143
rect 1008 -162 1024 -145
rect 1026 -162 1031 -137
rect 1033 -146 1038 -137
rect 1045 -138 1048 -136
rect 1050 -138 1054 -136
rect 1045 -146 1054 -138
rect 1033 -155 1041 -146
rect 1033 -157 1036 -155
rect 1038 -157 1041 -155
rect 1033 -159 1041 -157
rect 1043 -159 1054 -146
rect 1056 -146 1061 -134
rect 1070 -141 1075 -134
rect 1068 -143 1075 -141
rect 1068 -145 1070 -143
rect 1072 -145 1075 -143
rect 1056 -148 1063 -146
rect 1068 -147 1075 -145
rect 1056 -150 1059 -148
rect 1061 -150 1063 -148
rect 1056 -155 1063 -150
rect 1070 -155 1075 -147
rect 1077 -155 1082 -134
rect 1084 -136 1093 -134
rect 1084 -138 1089 -136
rect 1091 -138 1093 -136
rect 1084 -144 1093 -138
rect 1116 -143 1123 -141
rect 1084 -155 1095 -144
rect 1056 -157 1059 -155
rect 1061 -157 1063 -155
rect 1056 -159 1063 -157
rect 1033 -162 1038 -159
rect 1087 -162 1095 -155
rect 1097 -146 1104 -144
rect 1097 -148 1100 -146
rect 1102 -148 1104 -146
rect 1097 -153 1104 -148
rect 1097 -155 1100 -153
rect 1102 -155 1104 -153
rect 1116 -145 1118 -143
rect 1120 -145 1123 -143
rect 1116 -154 1123 -145
rect 1125 -143 1133 -141
rect 1125 -145 1128 -143
rect 1130 -145 1133 -143
rect 1125 -150 1133 -145
rect 1125 -152 1128 -150
rect 1130 -152 1133 -150
rect 1125 -154 1133 -152
rect 1135 -143 1141 -141
rect 1135 -145 1143 -143
rect 1135 -147 1138 -145
rect 1140 -147 1143 -145
rect 1135 -154 1143 -147
rect 1097 -157 1104 -155
rect 1097 -162 1102 -157
rect 1137 -161 1143 -154
rect 1145 -148 1150 -143
rect 1158 -146 1163 -134
rect 1156 -148 1163 -146
rect 1145 -150 1152 -148
rect 1145 -152 1148 -150
rect 1150 -152 1152 -150
rect 1145 -157 1152 -152
rect 1145 -159 1148 -157
rect 1150 -159 1152 -157
rect 1156 -150 1158 -148
rect 1160 -150 1163 -148
rect 1156 -155 1163 -150
rect 1156 -157 1158 -155
rect 1160 -157 1163 -155
rect 1156 -159 1163 -157
rect 1165 -136 1174 -134
rect 1165 -138 1169 -136
rect 1171 -138 1174 -136
rect 1197 -136 1211 -134
rect 1197 -137 1204 -136
rect 1165 -146 1174 -138
rect 1181 -146 1186 -137
rect 1165 -159 1176 -146
rect 1178 -155 1186 -146
rect 1178 -157 1181 -155
rect 1183 -157 1186 -155
rect 1178 -159 1186 -157
rect 1145 -161 1152 -159
rect 1181 -162 1186 -159
rect 1188 -162 1193 -137
rect 1195 -138 1204 -137
rect 1206 -138 1211 -136
rect 1195 -143 1211 -138
rect 1195 -145 1204 -143
rect 1206 -145 1211 -143
rect 1195 -162 1211 -145
rect 1213 -144 1221 -134
rect 1213 -146 1216 -144
rect 1218 -146 1221 -144
rect 1213 -151 1221 -146
rect 1213 -153 1216 -151
rect 1218 -153 1221 -151
rect 1213 -162 1221 -153
rect 1223 -136 1231 -134
rect 1223 -138 1226 -136
rect 1228 -138 1231 -136
rect 1223 -143 1231 -138
rect 1223 -145 1226 -143
rect 1228 -145 1231 -143
rect 1223 -162 1231 -145
rect 1233 -149 1238 -134
rect 1248 -149 1253 -134
rect 1233 -151 1240 -149
rect 1233 -153 1236 -151
rect 1238 -153 1240 -151
rect 1233 -158 1240 -153
rect 1233 -160 1236 -158
rect 1238 -160 1240 -158
rect 1233 -162 1240 -160
rect 1246 -151 1253 -149
rect 1246 -153 1248 -151
rect 1250 -153 1253 -151
rect 1246 -158 1253 -153
rect 1246 -160 1248 -158
rect 1250 -160 1253 -158
rect 1246 -162 1253 -160
rect 1255 -136 1263 -134
rect 1255 -138 1258 -136
rect 1260 -138 1263 -136
rect 1255 -143 1263 -138
rect 1255 -145 1258 -143
rect 1260 -145 1263 -143
rect 1255 -162 1263 -145
rect 1265 -144 1273 -134
rect 1265 -146 1268 -144
rect 1270 -146 1273 -144
rect 1265 -151 1273 -146
rect 1265 -153 1268 -151
rect 1270 -153 1273 -151
rect 1265 -162 1273 -153
rect 1275 -136 1289 -134
rect 1275 -138 1280 -136
rect 1282 -137 1289 -136
rect 1312 -136 1321 -134
rect 1282 -138 1291 -137
rect 1275 -143 1291 -138
rect 1275 -145 1280 -143
rect 1282 -145 1291 -143
rect 1275 -162 1291 -145
rect 1293 -162 1298 -137
rect 1300 -146 1305 -137
rect 1312 -138 1315 -136
rect 1317 -138 1321 -136
rect 1312 -146 1321 -138
rect 1300 -155 1308 -146
rect 1300 -157 1303 -155
rect 1305 -157 1308 -155
rect 1300 -159 1308 -157
rect 1310 -159 1321 -146
rect 1323 -146 1328 -134
rect 1337 -141 1342 -134
rect 1335 -143 1342 -141
rect 1335 -145 1337 -143
rect 1339 -145 1342 -143
rect 1323 -148 1330 -146
rect 1335 -147 1342 -145
rect 1323 -150 1326 -148
rect 1328 -150 1330 -148
rect 1323 -155 1330 -150
rect 1337 -155 1342 -147
rect 1344 -155 1349 -134
rect 1351 -136 1360 -134
rect 1351 -138 1356 -136
rect 1358 -138 1360 -136
rect 1351 -144 1360 -138
rect 1383 -143 1390 -141
rect 1351 -155 1362 -144
rect 1323 -157 1326 -155
rect 1328 -157 1330 -155
rect 1323 -159 1330 -157
rect 1300 -162 1305 -159
rect 1354 -162 1362 -155
rect 1364 -146 1371 -144
rect 1364 -148 1367 -146
rect 1369 -148 1371 -146
rect 1364 -153 1371 -148
rect 1364 -155 1367 -153
rect 1369 -155 1371 -153
rect 1383 -145 1385 -143
rect 1387 -145 1390 -143
rect 1383 -154 1390 -145
rect 1392 -143 1400 -141
rect 1392 -145 1395 -143
rect 1397 -145 1400 -143
rect 1392 -150 1400 -145
rect 1392 -152 1395 -150
rect 1397 -152 1400 -150
rect 1392 -154 1400 -152
rect 1402 -143 1408 -141
rect 1402 -145 1410 -143
rect 1402 -147 1405 -145
rect 1407 -147 1410 -145
rect 1402 -154 1410 -147
rect 1364 -157 1371 -155
rect 1364 -162 1369 -157
rect 1404 -161 1410 -154
rect 1412 -148 1417 -143
rect 1425 -146 1430 -134
rect 1423 -148 1430 -146
rect 1412 -150 1419 -148
rect 1412 -152 1415 -150
rect 1417 -152 1419 -150
rect 1412 -157 1419 -152
rect 1412 -159 1415 -157
rect 1417 -159 1419 -157
rect 1423 -150 1425 -148
rect 1427 -150 1430 -148
rect 1423 -155 1430 -150
rect 1423 -157 1425 -155
rect 1427 -157 1430 -155
rect 1423 -159 1430 -157
rect 1432 -136 1441 -134
rect 1432 -138 1436 -136
rect 1438 -138 1441 -136
rect 1464 -136 1478 -134
rect 1464 -137 1471 -136
rect 1432 -146 1441 -138
rect 1448 -146 1453 -137
rect 1432 -159 1443 -146
rect 1445 -155 1453 -146
rect 1445 -157 1448 -155
rect 1450 -157 1453 -155
rect 1445 -159 1453 -157
rect 1412 -161 1419 -159
rect 1448 -162 1453 -159
rect 1455 -162 1460 -137
rect 1462 -138 1471 -137
rect 1473 -138 1478 -136
rect 1462 -143 1478 -138
rect 1462 -145 1471 -143
rect 1473 -145 1478 -143
rect 1462 -162 1478 -145
rect 1480 -144 1488 -134
rect 1480 -146 1483 -144
rect 1485 -146 1488 -144
rect 1480 -151 1488 -146
rect 1480 -153 1483 -151
rect 1485 -153 1488 -151
rect 1480 -162 1488 -153
rect 1490 -136 1498 -134
rect 1490 -138 1493 -136
rect 1495 -138 1498 -136
rect 1490 -143 1498 -138
rect 1490 -145 1493 -143
rect 1495 -145 1498 -143
rect 1490 -162 1498 -145
rect 1500 -149 1505 -134
rect 1515 -149 1520 -134
rect 1500 -151 1507 -149
rect 1500 -153 1503 -151
rect 1505 -153 1507 -151
rect 1500 -158 1507 -153
rect 1500 -160 1503 -158
rect 1505 -160 1507 -158
rect 1500 -162 1507 -160
rect 1513 -151 1520 -149
rect 1513 -153 1515 -151
rect 1517 -153 1520 -151
rect 1513 -158 1520 -153
rect 1513 -160 1515 -158
rect 1517 -160 1520 -158
rect 1513 -162 1520 -160
rect 1522 -136 1530 -134
rect 1522 -138 1525 -136
rect 1527 -138 1530 -136
rect 1522 -143 1530 -138
rect 1522 -145 1525 -143
rect 1527 -145 1530 -143
rect 1522 -162 1530 -145
rect 1532 -144 1540 -134
rect 1532 -146 1535 -144
rect 1537 -146 1540 -144
rect 1532 -151 1540 -146
rect 1532 -153 1535 -151
rect 1537 -153 1540 -151
rect 1532 -162 1540 -153
rect 1542 -136 1556 -134
rect 1542 -138 1547 -136
rect 1549 -137 1556 -136
rect 1579 -136 1588 -134
rect 1549 -138 1558 -137
rect 1542 -143 1558 -138
rect 1542 -145 1547 -143
rect 1549 -145 1558 -143
rect 1542 -162 1558 -145
rect 1560 -162 1565 -137
rect 1567 -146 1572 -137
rect 1579 -138 1582 -136
rect 1584 -138 1588 -136
rect 1579 -146 1588 -138
rect 1567 -155 1575 -146
rect 1567 -157 1570 -155
rect 1572 -157 1575 -155
rect 1567 -159 1575 -157
rect 1577 -159 1588 -146
rect 1590 -146 1595 -134
rect 1604 -141 1609 -134
rect 1602 -143 1609 -141
rect 1602 -145 1604 -143
rect 1606 -145 1609 -143
rect 1590 -148 1597 -146
rect 1602 -147 1609 -145
rect 1590 -150 1593 -148
rect 1595 -150 1597 -148
rect 1590 -155 1597 -150
rect 1604 -155 1609 -147
rect 1611 -155 1616 -134
rect 1618 -136 1627 -134
rect 1618 -138 1623 -136
rect 1625 -138 1627 -136
rect 1618 -144 1627 -138
rect 1650 -143 1657 -141
rect 1618 -155 1629 -144
rect 1590 -157 1593 -155
rect 1595 -157 1597 -155
rect 1590 -159 1597 -157
rect 1567 -162 1572 -159
rect 1621 -162 1629 -155
rect 1631 -146 1638 -144
rect 1631 -148 1634 -146
rect 1636 -148 1638 -146
rect 1631 -153 1638 -148
rect 1631 -155 1634 -153
rect 1636 -155 1638 -153
rect 1650 -145 1652 -143
rect 1654 -145 1657 -143
rect 1650 -154 1657 -145
rect 1659 -143 1667 -141
rect 1659 -145 1662 -143
rect 1664 -145 1667 -143
rect 1659 -150 1667 -145
rect 1659 -152 1662 -150
rect 1664 -152 1667 -150
rect 1659 -154 1667 -152
rect 1669 -143 1675 -141
rect 1669 -145 1677 -143
rect 1669 -147 1672 -145
rect 1674 -147 1677 -145
rect 1669 -154 1677 -147
rect 1631 -157 1638 -155
rect 1631 -162 1636 -157
rect 1671 -161 1677 -154
rect 1679 -148 1684 -143
rect 1692 -146 1697 -134
rect 1690 -148 1697 -146
rect 1679 -150 1686 -148
rect 1679 -152 1682 -150
rect 1684 -152 1686 -150
rect 1679 -157 1686 -152
rect 1679 -159 1682 -157
rect 1684 -159 1686 -157
rect 1690 -150 1692 -148
rect 1694 -150 1697 -148
rect 1690 -155 1697 -150
rect 1690 -157 1692 -155
rect 1694 -157 1697 -155
rect 1690 -159 1697 -157
rect 1699 -136 1708 -134
rect 1699 -138 1703 -136
rect 1705 -138 1708 -136
rect 1731 -136 1745 -134
rect 1731 -137 1738 -136
rect 1699 -146 1708 -138
rect 1715 -146 1720 -137
rect 1699 -159 1710 -146
rect 1712 -155 1720 -146
rect 1712 -157 1715 -155
rect 1717 -157 1720 -155
rect 1712 -159 1720 -157
rect 1679 -161 1686 -159
rect 1715 -162 1720 -159
rect 1722 -162 1727 -137
rect 1729 -138 1738 -137
rect 1740 -138 1745 -136
rect 1729 -143 1745 -138
rect 1729 -145 1738 -143
rect 1740 -145 1745 -143
rect 1729 -162 1745 -145
rect 1747 -144 1755 -134
rect 1747 -146 1750 -144
rect 1752 -146 1755 -144
rect 1747 -151 1755 -146
rect 1747 -153 1750 -151
rect 1752 -153 1755 -151
rect 1747 -162 1755 -153
rect 1757 -136 1765 -134
rect 1757 -138 1760 -136
rect 1762 -138 1765 -136
rect 1757 -143 1765 -138
rect 1757 -145 1760 -143
rect 1762 -145 1765 -143
rect 1757 -162 1765 -145
rect 1767 -149 1772 -134
rect 1782 -149 1787 -134
rect 1767 -151 1774 -149
rect 1767 -153 1770 -151
rect 1772 -153 1774 -151
rect 1767 -158 1774 -153
rect 1767 -160 1770 -158
rect 1772 -160 1774 -158
rect 1767 -162 1774 -160
rect 1780 -151 1787 -149
rect 1780 -153 1782 -151
rect 1784 -153 1787 -151
rect 1780 -158 1787 -153
rect 1780 -160 1782 -158
rect 1784 -160 1787 -158
rect 1780 -162 1787 -160
rect 1789 -136 1797 -134
rect 1789 -138 1792 -136
rect 1794 -138 1797 -136
rect 1789 -143 1797 -138
rect 1789 -145 1792 -143
rect 1794 -145 1797 -143
rect 1789 -162 1797 -145
rect 1799 -144 1807 -134
rect 1799 -146 1802 -144
rect 1804 -146 1807 -144
rect 1799 -151 1807 -146
rect 1799 -153 1802 -151
rect 1804 -153 1807 -151
rect 1799 -162 1807 -153
rect 1809 -136 1823 -134
rect 1809 -138 1814 -136
rect 1816 -137 1823 -136
rect 1846 -136 1855 -134
rect 1816 -138 1825 -137
rect 1809 -143 1825 -138
rect 1809 -145 1814 -143
rect 1816 -145 1825 -143
rect 1809 -162 1825 -145
rect 1827 -162 1832 -137
rect 1834 -146 1839 -137
rect 1846 -138 1849 -136
rect 1851 -138 1855 -136
rect 1846 -146 1855 -138
rect 1834 -155 1842 -146
rect 1834 -157 1837 -155
rect 1839 -157 1842 -155
rect 1834 -159 1842 -157
rect 1844 -159 1855 -146
rect 1857 -146 1862 -134
rect 1871 -141 1876 -134
rect 1869 -143 1876 -141
rect 1869 -145 1871 -143
rect 1873 -145 1876 -143
rect 1857 -148 1864 -146
rect 1869 -147 1876 -145
rect 1857 -150 1860 -148
rect 1862 -150 1864 -148
rect 1857 -155 1864 -150
rect 1871 -155 1876 -147
rect 1878 -155 1883 -134
rect 1885 -136 1894 -134
rect 1885 -138 1890 -136
rect 1892 -138 1894 -136
rect 1885 -144 1894 -138
rect 1885 -155 1896 -144
rect 1857 -157 1860 -155
rect 1862 -157 1864 -155
rect 1857 -159 1864 -157
rect 1834 -162 1839 -159
rect 1888 -162 1896 -155
rect 1898 -146 1905 -144
rect 1898 -148 1901 -146
rect 1903 -148 1905 -146
rect 1898 -153 1905 -148
rect 1898 -155 1901 -153
rect 1903 -155 1905 -153
rect 1922 -155 1927 -134
rect 1898 -157 1905 -155
rect 1920 -157 1927 -155
rect 1898 -162 1903 -157
rect 1920 -159 1922 -157
rect 1924 -159 1927 -157
rect 1920 -161 1927 -159
rect 1929 -136 1941 -134
rect 1929 -138 1932 -136
rect 1934 -138 1941 -136
rect 1929 -143 1941 -138
rect 1958 -143 1963 -134
rect 1929 -145 1932 -143
rect 1934 -145 1943 -143
rect 1929 -161 1943 -145
rect 1945 -150 1953 -143
rect 1945 -152 1948 -150
rect 1950 -152 1953 -150
rect 1945 -157 1953 -152
rect 1945 -159 1948 -157
rect 1950 -159 1953 -157
rect 1945 -161 1953 -159
rect 1955 -150 1963 -143
rect 1955 -152 1958 -150
rect 1960 -152 1963 -150
rect 1955 -161 1963 -152
rect 1965 -140 1970 -134
rect 1965 -142 1972 -140
rect 1965 -144 1968 -142
rect 1970 -144 1972 -142
rect 1965 -146 1972 -144
rect 1978 -146 1983 -134
rect 1965 -161 1970 -146
rect 1976 -148 1983 -146
rect 1976 -150 1978 -148
rect 1980 -150 1983 -148
rect 1976 -155 1983 -150
rect 1976 -157 1978 -155
rect 1980 -157 1983 -155
rect 1976 -159 1983 -157
rect 1985 -136 1994 -134
rect 1985 -138 1989 -136
rect 1991 -138 1994 -136
rect 2017 -136 2031 -134
rect 2017 -137 2024 -136
rect 1985 -146 1994 -138
rect 2001 -146 2006 -137
rect 1985 -159 1996 -146
rect 1998 -155 2006 -146
rect 1998 -157 2001 -155
rect 2003 -157 2006 -155
rect 1998 -159 2006 -157
rect 2001 -162 2006 -159
rect 2008 -162 2013 -137
rect 2015 -138 2024 -137
rect 2026 -138 2031 -136
rect 2015 -143 2031 -138
rect 2015 -145 2024 -143
rect 2026 -145 2031 -143
rect 2015 -162 2031 -145
rect 2033 -144 2041 -134
rect 2033 -146 2036 -144
rect 2038 -146 2041 -144
rect 2033 -151 2041 -146
rect 2033 -153 2036 -151
rect 2038 -153 2041 -151
rect 2033 -162 2041 -153
rect 2043 -136 2051 -134
rect 2043 -138 2046 -136
rect 2048 -138 2051 -136
rect 2043 -143 2051 -138
rect 2043 -145 2046 -143
rect 2048 -145 2051 -143
rect 2043 -162 2051 -145
rect 2053 -149 2058 -134
rect 2068 -149 2073 -134
rect 2053 -151 2060 -149
rect 2053 -153 2056 -151
rect 2058 -153 2060 -151
rect 2053 -158 2060 -153
rect 2053 -160 2056 -158
rect 2058 -160 2060 -158
rect 2053 -162 2060 -160
rect 2066 -151 2073 -149
rect 2066 -153 2068 -151
rect 2070 -153 2073 -151
rect 2066 -158 2073 -153
rect 2066 -160 2068 -158
rect 2070 -160 2073 -158
rect 2066 -162 2073 -160
rect 2075 -136 2083 -134
rect 2075 -138 2078 -136
rect 2080 -138 2083 -136
rect 2075 -143 2083 -138
rect 2075 -145 2078 -143
rect 2080 -145 2083 -143
rect 2075 -162 2083 -145
rect 2085 -144 2093 -134
rect 2085 -146 2088 -144
rect 2090 -146 2093 -144
rect 2085 -151 2093 -146
rect 2085 -153 2088 -151
rect 2090 -153 2093 -151
rect 2085 -162 2093 -153
rect 2095 -136 2109 -134
rect 2095 -138 2100 -136
rect 2102 -137 2109 -136
rect 2132 -136 2141 -134
rect 2102 -138 2111 -137
rect 2095 -143 2111 -138
rect 2095 -145 2100 -143
rect 2102 -145 2111 -143
rect 2095 -162 2111 -145
rect 2113 -162 2118 -137
rect 2120 -146 2125 -137
rect 2132 -138 2135 -136
rect 2137 -138 2141 -136
rect 2132 -146 2141 -138
rect 2120 -155 2128 -146
rect 2120 -157 2123 -155
rect 2125 -157 2128 -155
rect 2120 -159 2128 -157
rect 2130 -159 2141 -146
rect 2143 -146 2148 -134
rect 2157 -141 2162 -134
rect 2155 -143 2162 -141
rect 2155 -145 2157 -143
rect 2159 -145 2162 -143
rect 2143 -148 2150 -146
rect 2155 -147 2162 -145
rect 2143 -150 2146 -148
rect 2148 -150 2150 -148
rect 2143 -155 2150 -150
rect 2157 -155 2162 -147
rect 2164 -155 2169 -134
rect 2171 -136 2180 -134
rect 2171 -138 2176 -136
rect 2178 -138 2180 -136
rect 2209 -136 2216 -134
rect 2171 -144 2180 -138
rect 2209 -138 2211 -136
rect 2213 -138 2216 -136
rect 2171 -155 2182 -144
rect 2143 -157 2146 -155
rect 2148 -157 2150 -155
rect 2143 -159 2150 -157
rect 2120 -162 2125 -159
rect 2174 -162 2182 -155
rect 2184 -146 2191 -144
rect 2184 -148 2187 -146
rect 2189 -148 2191 -146
rect 2184 -153 2191 -148
rect 2209 -146 2216 -138
rect 2184 -155 2187 -153
rect 2189 -155 2191 -153
rect 2210 -150 2216 -146
rect 2218 -150 2223 -134
rect 2225 -146 2233 -134
rect 2225 -148 2228 -146
rect 2230 -148 2233 -146
rect 2225 -150 2233 -148
rect 2235 -150 2240 -134
rect 2242 -136 2250 -134
rect 2242 -138 2245 -136
rect 2247 -138 2250 -136
rect 2242 -150 2250 -138
rect 2210 -154 2214 -150
rect 2184 -157 2191 -155
rect 2201 -156 2206 -154
rect 2184 -162 2189 -157
rect 2199 -158 2206 -156
rect 2199 -160 2201 -158
rect 2203 -160 2206 -158
rect 2199 -162 2206 -160
rect 2208 -162 2214 -154
rect 2245 -152 2250 -150
rect 2252 -141 2257 -134
rect 2277 -136 2284 -134
rect 2277 -138 2279 -136
rect 2281 -138 2284 -136
rect 2252 -143 2259 -141
rect 2252 -145 2255 -143
rect 2257 -145 2259 -143
rect 2252 -147 2259 -145
rect 2277 -146 2284 -138
rect 2252 -152 2257 -147
rect 2278 -150 2284 -146
rect 2286 -150 2291 -134
rect 2293 -146 2301 -134
rect 2293 -148 2296 -146
rect 2298 -148 2301 -146
rect 2293 -150 2301 -148
rect 2303 -150 2308 -134
rect 2310 -136 2318 -134
rect 2310 -138 2313 -136
rect 2315 -138 2318 -136
rect 2310 -150 2318 -138
rect 2278 -154 2282 -150
rect 2269 -156 2274 -154
rect 2267 -158 2274 -156
rect 2267 -160 2269 -158
rect 2271 -160 2274 -158
rect 2267 -162 2274 -160
rect 2276 -162 2282 -154
rect 2313 -152 2318 -150
rect 2320 -141 2325 -134
rect 2320 -143 2327 -141
rect 2320 -145 2323 -143
rect 2325 -145 2327 -143
rect 2320 -147 2327 -145
rect 2320 -152 2325 -147
rect 29 -246 35 -239
rect 8 -255 15 -246
rect 8 -257 10 -255
rect 12 -257 15 -255
rect 8 -259 15 -257
rect 17 -248 25 -246
rect 17 -250 20 -248
rect 22 -250 25 -248
rect 17 -255 25 -250
rect 17 -257 20 -255
rect 22 -257 25 -255
rect 17 -259 25 -257
rect 27 -253 35 -246
rect 27 -255 30 -253
rect 32 -255 35 -253
rect 27 -257 35 -255
rect 37 -241 44 -239
rect 37 -243 40 -241
rect 42 -243 44 -241
rect 37 -248 44 -243
rect 69 -246 75 -239
rect 37 -250 40 -248
rect 42 -250 44 -248
rect 37 -252 44 -250
rect 37 -257 42 -252
rect 48 -255 55 -246
rect 48 -257 50 -255
rect 52 -257 55 -255
rect 27 -259 33 -257
rect 48 -259 55 -257
rect 57 -248 65 -246
rect 57 -250 60 -248
rect 62 -250 65 -248
rect 57 -255 65 -250
rect 57 -257 60 -255
rect 62 -257 65 -255
rect 57 -259 65 -257
rect 67 -253 75 -246
rect 67 -255 70 -253
rect 72 -255 75 -253
rect 67 -257 75 -255
rect 77 -241 84 -239
rect 113 -241 118 -238
rect 77 -243 80 -241
rect 82 -243 84 -241
rect 77 -248 84 -243
rect 77 -250 80 -248
rect 82 -250 84 -248
rect 77 -252 84 -250
rect 88 -243 95 -241
rect 88 -245 90 -243
rect 92 -245 95 -243
rect 88 -250 95 -245
rect 88 -252 90 -250
rect 92 -252 95 -250
rect 77 -257 82 -252
rect 88 -254 95 -252
rect 67 -259 73 -257
rect 90 -266 95 -254
rect 97 -254 108 -241
rect 110 -243 118 -241
rect 110 -245 113 -243
rect 115 -245 118 -243
rect 110 -254 118 -245
rect 97 -262 106 -254
rect 97 -264 101 -262
rect 103 -264 106 -262
rect 113 -263 118 -254
rect 120 -263 125 -238
rect 127 -255 143 -238
rect 127 -257 136 -255
rect 138 -257 143 -255
rect 127 -262 143 -257
rect 127 -263 136 -262
rect 97 -266 106 -264
rect 129 -264 136 -263
rect 138 -264 143 -262
rect 129 -266 143 -264
rect 145 -247 153 -238
rect 145 -249 148 -247
rect 150 -249 153 -247
rect 145 -254 153 -249
rect 145 -256 148 -254
rect 150 -256 153 -254
rect 145 -266 153 -256
rect 155 -255 163 -238
rect 155 -257 158 -255
rect 160 -257 163 -255
rect 155 -262 163 -257
rect 155 -264 158 -262
rect 160 -264 163 -262
rect 155 -266 163 -264
rect 165 -240 172 -238
rect 165 -242 168 -240
rect 170 -242 172 -240
rect 165 -247 172 -242
rect 165 -249 168 -247
rect 170 -249 172 -247
rect 165 -251 172 -249
rect 178 -240 185 -238
rect 178 -242 180 -240
rect 182 -242 185 -240
rect 178 -247 185 -242
rect 178 -249 180 -247
rect 182 -249 185 -247
rect 178 -251 185 -249
rect 165 -266 170 -251
rect 180 -266 185 -251
rect 187 -255 195 -238
rect 187 -257 190 -255
rect 192 -257 195 -255
rect 187 -262 195 -257
rect 187 -264 190 -262
rect 192 -264 195 -262
rect 187 -266 195 -264
rect 197 -247 205 -238
rect 197 -249 200 -247
rect 202 -249 205 -247
rect 197 -254 205 -249
rect 197 -256 200 -254
rect 202 -256 205 -254
rect 197 -266 205 -256
rect 207 -255 223 -238
rect 207 -257 212 -255
rect 214 -257 223 -255
rect 207 -262 223 -257
rect 207 -264 212 -262
rect 214 -263 223 -262
rect 225 -263 230 -238
rect 232 -241 237 -238
rect 232 -243 240 -241
rect 232 -245 235 -243
rect 237 -245 240 -243
rect 232 -254 240 -245
rect 242 -254 253 -241
rect 232 -263 237 -254
rect 244 -262 253 -254
rect 214 -264 221 -263
rect 207 -266 221 -264
rect 244 -264 247 -262
rect 249 -264 253 -262
rect 244 -266 253 -264
rect 255 -243 262 -241
rect 255 -245 258 -243
rect 260 -245 262 -243
rect 286 -245 294 -238
rect 255 -250 262 -245
rect 255 -252 258 -250
rect 260 -252 262 -250
rect 255 -254 262 -252
rect 269 -253 274 -245
rect 255 -266 260 -254
rect 267 -255 274 -253
rect 267 -257 269 -255
rect 271 -257 274 -255
rect 267 -259 274 -257
rect 269 -266 274 -259
rect 276 -266 281 -245
rect 283 -256 294 -245
rect 296 -243 301 -238
rect 296 -245 303 -243
rect 296 -247 299 -245
rect 301 -247 303 -245
rect 336 -246 342 -239
rect 296 -252 303 -247
rect 296 -254 299 -252
rect 301 -254 303 -252
rect 296 -256 303 -254
rect 315 -255 322 -246
rect 283 -262 292 -256
rect 315 -257 317 -255
rect 319 -257 322 -255
rect 315 -259 322 -257
rect 324 -248 332 -246
rect 324 -250 327 -248
rect 329 -250 332 -248
rect 324 -255 332 -250
rect 324 -257 327 -255
rect 329 -257 332 -255
rect 324 -259 332 -257
rect 334 -253 342 -246
rect 334 -255 337 -253
rect 339 -255 342 -253
rect 334 -257 342 -255
rect 344 -241 351 -239
rect 380 -241 385 -238
rect 344 -243 347 -241
rect 349 -243 351 -241
rect 344 -248 351 -243
rect 344 -250 347 -248
rect 349 -250 351 -248
rect 344 -252 351 -250
rect 355 -243 362 -241
rect 355 -245 357 -243
rect 359 -245 362 -243
rect 355 -250 362 -245
rect 355 -252 357 -250
rect 359 -252 362 -250
rect 344 -257 349 -252
rect 355 -254 362 -252
rect 334 -259 340 -257
rect 283 -264 288 -262
rect 290 -264 292 -262
rect 283 -266 292 -264
rect 357 -266 362 -254
rect 364 -254 375 -241
rect 377 -243 385 -241
rect 377 -245 380 -243
rect 382 -245 385 -243
rect 377 -254 385 -245
rect 364 -262 373 -254
rect 364 -264 368 -262
rect 370 -264 373 -262
rect 380 -263 385 -254
rect 387 -263 392 -238
rect 394 -255 410 -238
rect 394 -257 403 -255
rect 405 -257 410 -255
rect 394 -262 410 -257
rect 394 -263 403 -262
rect 364 -266 373 -264
rect 396 -264 403 -263
rect 405 -264 410 -262
rect 396 -266 410 -264
rect 412 -247 420 -238
rect 412 -249 415 -247
rect 417 -249 420 -247
rect 412 -254 420 -249
rect 412 -256 415 -254
rect 417 -256 420 -254
rect 412 -266 420 -256
rect 422 -255 430 -238
rect 422 -257 425 -255
rect 427 -257 430 -255
rect 422 -262 430 -257
rect 422 -264 425 -262
rect 427 -264 430 -262
rect 422 -266 430 -264
rect 432 -240 439 -238
rect 432 -242 435 -240
rect 437 -242 439 -240
rect 432 -247 439 -242
rect 432 -249 435 -247
rect 437 -249 439 -247
rect 432 -251 439 -249
rect 445 -240 452 -238
rect 445 -242 447 -240
rect 449 -242 452 -240
rect 445 -247 452 -242
rect 445 -249 447 -247
rect 449 -249 452 -247
rect 445 -251 452 -249
rect 432 -266 437 -251
rect 447 -266 452 -251
rect 454 -255 462 -238
rect 454 -257 457 -255
rect 459 -257 462 -255
rect 454 -262 462 -257
rect 454 -264 457 -262
rect 459 -264 462 -262
rect 454 -266 462 -264
rect 464 -247 472 -238
rect 464 -249 467 -247
rect 469 -249 472 -247
rect 464 -254 472 -249
rect 464 -256 467 -254
rect 469 -256 472 -254
rect 464 -266 472 -256
rect 474 -255 490 -238
rect 474 -257 479 -255
rect 481 -257 490 -255
rect 474 -262 490 -257
rect 474 -264 479 -262
rect 481 -263 490 -262
rect 492 -263 497 -238
rect 499 -241 504 -238
rect 499 -243 507 -241
rect 499 -245 502 -243
rect 504 -245 507 -243
rect 499 -254 507 -245
rect 509 -254 520 -241
rect 499 -263 504 -254
rect 511 -262 520 -254
rect 481 -264 488 -263
rect 474 -266 488 -264
rect 511 -264 514 -262
rect 516 -264 520 -262
rect 511 -266 520 -264
rect 522 -243 529 -241
rect 522 -245 525 -243
rect 527 -245 529 -243
rect 553 -245 561 -238
rect 522 -250 529 -245
rect 522 -252 525 -250
rect 527 -252 529 -250
rect 522 -254 529 -252
rect 536 -253 541 -245
rect 522 -266 527 -254
rect 534 -255 541 -253
rect 534 -257 536 -255
rect 538 -257 541 -255
rect 534 -259 541 -257
rect 536 -266 541 -259
rect 543 -266 548 -245
rect 550 -256 561 -245
rect 563 -243 568 -238
rect 563 -245 570 -243
rect 563 -247 566 -245
rect 568 -247 570 -245
rect 603 -246 609 -239
rect 563 -252 570 -247
rect 563 -254 566 -252
rect 568 -254 570 -252
rect 563 -256 570 -254
rect 582 -255 589 -246
rect 550 -262 559 -256
rect 582 -257 584 -255
rect 586 -257 589 -255
rect 582 -259 589 -257
rect 591 -248 599 -246
rect 591 -250 594 -248
rect 596 -250 599 -248
rect 591 -255 599 -250
rect 591 -257 594 -255
rect 596 -257 599 -255
rect 591 -259 599 -257
rect 601 -253 609 -246
rect 601 -255 604 -253
rect 606 -255 609 -253
rect 601 -257 609 -255
rect 611 -241 618 -239
rect 647 -241 652 -238
rect 611 -243 614 -241
rect 616 -243 618 -241
rect 611 -248 618 -243
rect 611 -250 614 -248
rect 616 -250 618 -248
rect 611 -252 618 -250
rect 622 -243 629 -241
rect 622 -245 624 -243
rect 626 -245 629 -243
rect 622 -250 629 -245
rect 622 -252 624 -250
rect 626 -252 629 -250
rect 611 -257 616 -252
rect 622 -254 629 -252
rect 601 -259 607 -257
rect 550 -264 555 -262
rect 557 -264 559 -262
rect 550 -266 559 -264
rect 624 -266 629 -254
rect 631 -254 642 -241
rect 644 -243 652 -241
rect 644 -245 647 -243
rect 649 -245 652 -243
rect 644 -254 652 -245
rect 631 -262 640 -254
rect 631 -264 635 -262
rect 637 -264 640 -262
rect 647 -263 652 -254
rect 654 -263 659 -238
rect 661 -255 677 -238
rect 661 -257 670 -255
rect 672 -257 677 -255
rect 661 -262 677 -257
rect 661 -263 670 -262
rect 631 -266 640 -264
rect 663 -264 670 -263
rect 672 -264 677 -262
rect 663 -266 677 -264
rect 679 -247 687 -238
rect 679 -249 682 -247
rect 684 -249 687 -247
rect 679 -254 687 -249
rect 679 -256 682 -254
rect 684 -256 687 -254
rect 679 -266 687 -256
rect 689 -255 697 -238
rect 689 -257 692 -255
rect 694 -257 697 -255
rect 689 -262 697 -257
rect 689 -264 692 -262
rect 694 -264 697 -262
rect 689 -266 697 -264
rect 699 -240 706 -238
rect 699 -242 702 -240
rect 704 -242 706 -240
rect 699 -247 706 -242
rect 699 -249 702 -247
rect 704 -249 706 -247
rect 699 -251 706 -249
rect 712 -240 719 -238
rect 712 -242 714 -240
rect 716 -242 719 -240
rect 712 -247 719 -242
rect 712 -249 714 -247
rect 716 -249 719 -247
rect 712 -251 719 -249
rect 699 -266 704 -251
rect 714 -266 719 -251
rect 721 -255 729 -238
rect 721 -257 724 -255
rect 726 -257 729 -255
rect 721 -262 729 -257
rect 721 -264 724 -262
rect 726 -264 729 -262
rect 721 -266 729 -264
rect 731 -247 739 -238
rect 731 -249 734 -247
rect 736 -249 739 -247
rect 731 -254 739 -249
rect 731 -256 734 -254
rect 736 -256 739 -254
rect 731 -266 739 -256
rect 741 -255 757 -238
rect 741 -257 746 -255
rect 748 -257 757 -255
rect 741 -262 757 -257
rect 741 -264 746 -262
rect 748 -263 757 -262
rect 759 -263 764 -238
rect 766 -241 771 -238
rect 766 -243 774 -241
rect 766 -245 769 -243
rect 771 -245 774 -243
rect 766 -254 774 -245
rect 776 -254 787 -241
rect 766 -263 771 -254
rect 778 -262 787 -254
rect 748 -264 755 -263
rect 741 -266 755 -264
rect 778 -264 781 -262
rect 783 -264 787 -262
rect 778 -266 787 -264
rect 789 -243 796 -241
rect 789 -245 792 -243
rect 794 -245 796 -243
rect 820 -245 828 -238
rect 789 -250 796 -245
rect 789 -252 792 -250
rect 794 -252 796 -250
rect 789 -254 796 -252
rect 803 -253 808 -245
rect 789 -266 794 -254
rect 801 -255 808 -253
rect 801 -257 803 -255
rect 805 -257 808 -255
rect 801 -259 808 -257
rect 803 -266 808 -259
rect 810 -266 815 -245
rect 817 -256 828 -245
rect 830 -243 835 -238
rect 830 -245 837 -243
rect 830 -247 833 -245
rect 835 -247 837 -245
rect 870 -246 876 -239
rect 830 -252 837 -247
rect 830 -254 833 -252
rect 835 -254 837 -252
rect 830 -256 837 -254
rect 849 -255 856 -246
rect 817 -262 826 -256
rect 849 -257 851 -255
rect 853 -257 856 -255
rect 849 -259 856 -257
rect 858 -248 866 -246
rect 858 -250 861 -248
rect 863 -250 866 -248
rect 858 -255 866 -250
rect 858 -257 861 -255
rect 863 -257 866 -255
rect 858 -259 866 -257
rect 868 -253 876 -246
rect 868 -255 871 -253
rect 873 -255 876 -253
rect 868 -257 876 -255
rect 878 -241 885 -239
rect 914 -241 919 -238
rect 878 -243 881 -241
rect 883 -243 885 -241
rect 878 -248 885 -243
rect 878 -250 881 -248
rect 883 -250 885 -248
rect 878 -252 885 -250
rect 889 -243 896 -241
rect 889 -245 891 -243
rect 893 -245 896 -243
rect 889 -250 896 -245
rect 889 -252 891 -250
rect 893 -252 896 -250
rect 878 -257 883 -252
rect 889 -254 896 -252
rect 868 -259 874 -257
rect 817 -264 822 -262
rect 824 -264 826 -262
rect 817 -266 826 -264
rect 891 -266 896 -254
rect 898 -254 909 -241
rect 911 -243 919 -241
rect 911 -245 914 -243
rect 916 -245 919 -243
rect 911 -254 919 -245
rect 898 -262 907 -254
rect 898 -264 902 -262
rect 904 -264 907 -262
rect 914 -263 919 -254
rect 921 -263 926 -238
rect 928 -255 944 -238
rect 928 -257 937 -255
rect 939 -257 944 -255
rect 928 -262 944 -257
rect 928 -263 937 -262
rect 898 -266 907 -264
rect 930 -264 937 -263
rect 939 -264 944 -262
rect 930 -266 944 -264
rect 946 -247 954 -238
rect 946 -249 949 -247
rect 951 -249 954 -247
rect 946 -254 954 -249
rect 946 -256 949 -254
rect 951 -256 954 -254
rect 946 -266 954 -256
rect 956 -255 964 -238
rect 956 -257 959 -255
rect 961 -257 964 -255
rect 956 -262 964 -257
rect 956 -264 959 -262
rect 961 -264 964 -262
rect 956 -266 964 -264
rect 966 -240 973 -238
rect 966 -242 969 -240
rect 971 -242 973 -240
rect 966 -247 973 -242
rect 966 -249 969 -247
rect 971 -249 973 -247
rect 966 -251 973 -249
rect 979 -240 986 -238
rect 979 -242 981 -240
rect 983 -242 986 -240
rect 979 -247 986 -242
rect 979 -249 981 -247
rect 983 -249 986 -247
rect 979 -251 986 -249
rect 966 -266 971 -251
rect 981 -266 986 -251
rect 988 -255 996 -238
rect 988 -257 991 -255
rect 993 -257 996 -255
rect 988 -262 996 -257
rect 988 -264 991 -262
rect 993 -264 996 -262
rect 988 -266 996 -264
rect 998 -247 1006 -238
rect 998 -249 1001 -247
rect 1003 -249 1006 -247
rect 998 -254 1006 -249
rect 998 -256 1001 -254
rect 1003 -256 1006 -254
rect 998 -266 1006 -256
rect 1008 -255 1024 -238
rect 1008 -257 1013 -255
rect 1015 -257 1024 -255
rect 1008 -262 1024 -257
rect 1008 -264 1013 -262
rect 1015 -263 1024 -262
rect 1026 -263 1031 -238
rect 1033 -241 1038 -238
rect 1033 -243 1041 -241
rect 1033 -245 1036 -243
rect 1038 -245 1041 -243
rect 1033 -254 1041 -245
rect 1043 -254 1054 -241
rect 1033 -263 1038 -254
rect 1045 -262 1054 -254
rect 1015 -264 1022 -263
rect 1008 -266 1022 -264
rect 1045 -264 1048 -262
rect 1050 -264 1054 -262
rect 1045 -266 1054 -264
rect 1056 -243 1063 -241
rect 1056 -245 1059 -243
rect 1061 -245 1063 -243
rect 1087 -245 1095 -238
rect 1056 -250 1063 -245
rect 1056 -252 1059 -250
rect 1061 -252 1063 -250
rect 1056 -254 1063 -252
rect 1070 -253 1075 -245
rect 1056 -266 1061 -254
rect 1068 -255 1075 -253
rect 1068 -257 1070 -255
rect 1072 -257 1075 -255
rect 1068 -259 1075 -257
rect 1070 -266 1075 -259
rect 1077 -266 1082 -245
rect 1084 -256 1095 -245
rect 1097 -243 1102 -238
rect 1097 -245 1104 -243
rect 1097 -247 1100 -245
rect 1102 -247 1104 -245
rect 1137 -246 1143 -239
rect 1097 -252 1104 -247
rect 1097 -254 1100 -252
rect 1102 -254 1104 -252
rect 1097 -256 1104 -254
rect 1116 -255 1123 -246
rect 1084 -262 1093 -256
rect 1116 -257 1118 -255
rect 1120 -257 1123 -255
rect 1116 -259 1123 -257
rect 1125 -248 1133 -246
rect 1125 -250 1128 -248
rect 1130 -250 1133 -248
rect 1125 -255 1133 -250
rect 1125 -257 1128 -255
rect 1130 -257 1133 -255
rect 1125 -259 1133 -257
rect 1135 -253 1143 -246
rect 1135 -255 1138 -253
rect 1140 -255 1143 -253
rect 1135 -257 1143 -255
rect 1145 -241 1152 -239
rect 1181 -241 1186 -238
rect 1145 -243 1148 -241
rect 1150 -243 1152 -241
rect 1145 -248 1152 -243
rect 1145 -250 1148 -248
rect 1150 -250 1152 -248
rect 1145 -252 1152 -250
rect 1156 -243 1163 -241
rect 1156 -245 1158 -243
rect 1160 -245 1163 -243
rect 1156 -250 1163 -245
rect 1156 -252 1158 -250
rect 1160 -252 1163 -250
rect 1145 -257 1150 -252
rect 1156 -254 1163 -252
rect 1135 -259 1141 -257
rect 1084 -264 1089 -262
rect 1091 -264 1093 -262
rect 1084 -266 1093 -264
rect 1158 -266 1163 -254
rect 1165 -254 1176 -241
rect 1178 -243 1186 -241
rect 1178 -245 1181 -243
rect 1183 -245 1186 -243
rect 1178 -254 1186 -245
rect 1165 -262 1174 -254
rect 1165 -264 1169 -262
rect 1171 -264 1174 -262
rect 1181 -263 1186 -254
rect 1188 -263 1193 -238
rect 1195 -255 1211 -238
rect 1195 -257 1204 -255
rect 1206 -257 1211 -255
rect 1195 -262 1211 -257
rect 1195 -263 1204 -262
rect 1165 -266 1174 -264
rect 1197 -264 1204 -263
rect 1206 -264 1211 -262
rect 1197 -266 1211 -264
rect 1213 -247 1221 -238
rect 1213 -249 1216 -247
rect 1218 -249 1221 -247
rect 1213 -254 1221 -249
rect 1213 -256 1216 -254
rect 1218 -256 1221 -254
rect 1213 -266 1221 -256
rect 1223 -255 1231 -238
rect 1223 -257 1226 -255
rect 1228 -257 1231 -255
rect 1223 -262 1231 -257
rect 1223 -264 1226 -262
rect 1228 -264 1231 -262
rect 1223 -266 1231 -264
rect 1233 -240 1240 -238
rect 1233 -242 1236 -240
rect 1238 -242 1240 -240
rect 1233 -247 1240 -242
rect 1233 -249 1236 -247
rect 1238 -249 1240 -247
rect 1233 -251 1240 -249
rect 1246 -240 1253 -238
rect 1246 -242 1248 -240
rect 1250 -242 1253 -240
rect 1246 -247 1253 -242
rect 1246 -249 1248 -247
rect 1250 -249 1253 -247
rect 1246 -251 1253 -249
rect 1233 -266 1238 -251
rect 1248 -266 1253 -251
rect 1255 -255 1263 -238
rect 1255 -257 1258 -255
rect 1260 -257 1263 -255
rect 1255 -262 1263 -257
rect 1255 -264 1258 -262
rect 1260 -264 1263 -262
rect 1255 -266 1263 -264
rect 1265 -247 1273 -238
rect 1265 -249 1268 -247
rect 1270 -249 1273 -247
rect 1265 -254 1273 -249
rect 1265 -256 1268 -254
rect 1270 -256 1273 -254
rect 1265 -266 1273 -256
rect 1275 -255 1291 -238
rect 1275 -257 1280 -255
rect 1282 -257 1291 -255
rect 1275 -262 1291 -257
rect 1275 -264 1280 -262
rect 1282 -263 1291 -262
rect 1293 -263 1298 -238
rect 1300 -241 1305 -238
rect 1300 -243 1308 -241
rect 1300 -245 1303 -243
rect 1305 -245 1308 -243
rect 1300 -254 1308 -245
rect 1310 -254 1321 -241
rect 1300 -263 1305 -254
rect 1312 -262 1321 -254
rect 1282 -264 1289 -263
rect 1275 -266 1289 -264
rect 1312 -264 1315 -262
rect 1317 -264 1321 -262
rect 1312 -266 1321 -264
rect 1323 -243 1330 -241
rect 1323 -245 1326 -243
rect 1328 -245 1330 -243
rect 1354 -245 1362 -238
rect 1323 -250 1330 -245
rect 1323 -252 1326 -250
rect 1328 -252 1330 -250
rect 1323 -254 1330 -252
rect 1337 -253 1342 -245
rect 1323 -266 1328 -254
rect 1335 -255 1342 -253
rect 1335 -257 1337 -255
rect 1339 -257 1342 -255
rect 1335 -259 1342 -257
rect 1337 -266 1342 -259
rect 1344 -266 1349 -245
rect 1351 -256 1362 -245
rect 1364 -243 1369 -238
rect 1364 -245 1371 -243
rect 1364 -247 1367 -245
rect 1369 -247 1371 -245
rect 1404 -246 1410 -239
rect 1364 -252 1371 -247
rect 1364 -254 1367 -252
rect 1369 -254 1371 -252
rect 1364 -256 1371 -254
rect 1383 -255 1390 -246
rect 1351 -262 1360 -256
rect 1383 -257 1385 -255
rect 1387 -257 1390 -255
rect 1383 -259 1390 -257
rect 1392 -248 1400 -246
rect 1392 -250 1395 -248
rect 1397 -250 1400 -248
rect 1392 -255 1400 -250
rect 1392 -257 1395 -255
rect 1397 -257 1400 -255
rect 1392 -259 1400 -257
rect 1402 -253 1410 -246
rect 1402 -255 1405 -253
rect 1407 -255 1410 -253
rect 1402 -257 1410 -255
rect 1412 -241 1419 -239
rect 1448 -241 1453 -238
rect 1412 -243 1415 -241
rect 1417 -243 1419 -241
rect 1412 -248 1419 -243
rect 1412 -250 1415 -248
rect 1417 -250 1419 -248
rect 1412 -252 1419 -250
rect 1423 -243 1430 -241
rect 1423 -245 1425 -243
rect 1427 -245 1430 -243
rect 1423 -250 1430 -245
rect 1423 -252 1425 -250
rect 1427 -252 1430 -250
rect 1412 -257 1417 -252
rect 1423 -254 1430 -252
rect 1402 -259 1408 -257
rect 1351 -264 1356 -262
rect 1358 -264 1360 -262
rect 1351 -266 1360 -264
rect 1425 -266 1430 -254
rect 1432 -254 1443 -241
rect 1445 -243 1453 -241
rect 1445 -245 1448 -243
rect 1450 -245 1453 -243
rect 1445 -254 1453 -245
rect 1432 -262 1441 -254
rect 1432 -264 1436 -262
rect 1438 -264 1441 -262
rect 1448 -263 1453 -254
rect 1455 -263 1460 -238
rect 1462 -255 1478 -238
rect 1462 -257 1471 -255
rect 1473 -257 1478 -255
rect 1462 -262 1478 -257
rect 1462 -263 1471 -262
rect 1432 -266 1441 -264
rect 1464 -264 1471 -263
rect 1473 -264 1478 -262
rect 1464 -266 1478 -264
rect 1480 -247 1488 -238
rect 1480 -249 1483 -247
rect 1485 -249 1488 -247
rect 1480 -254 1488 -249
rect 1480 -256 1483 -254
rect 1485 -256 1488 -254
rect 1480 -266 1488 -256
rect 1490 -255 1498 -238
rect 1490 -257 1493 -255
rect 1495 -257 1498 -255
rect 1490 -262 1498 -257
rect 1490 -264 1493 -262
rect 1495 -264 1498 -262
rect 1490 -266 1498 -264
rect 1500 -240 1507 -238
rect 1500 -242 1503 -240
rect 1505 -242 1507 -240
rect 1500 -247 1507 -242
rect 1500 -249 1503 -247
rect 1505 -249 1507 -247
rect 1500 -251 1507 -249
rect 1513 -240 1520 -238
rect 1513 -242 1515 -240
rect 1517 -242 1520 -240
rect 1513 -247 1520 -242
rect 1513 -249 1515 -247
rect 1517 -249 1520 -247
rect 1513 -251 1520 -249
rect 1500 -266 1505 -251
rect 1515 -266 1520 -251
rect 1522 -255 1530 -238
rect 1522 -257 1525 -255
rect 1527 -257 1530 -255
rect 1522 -262 1530 -257
rect 1522 -264 1525 -262
rect 1527 -264 1530 -262
rect 1522 -266 1530 -264
rect 1532 -247 1540 -238
rect 1532 -249 1535 -247
rect 1537 -249 1540 -247
rect 1532 -254 1540 -249
rect 1532 -256 1535 -254
rect 1537 -256 1540 -254
rect 1532 -266 1540 -256
rect 1542 -255 1558 -238
rect 1542 -257 1547 -255
rect 1549 -257 1558 -255
rect 1542 -262 1558 -257
rect 1542 -264 1547 -262
rect 1549 -263 1558 -262
rect 1560 -263 1565 -238
rect 1567 -241 1572 -238
rect 1567 -243 1575 -241
rect 1567 -245 1570 -243
rect 1572 -245 1575 -243
rect 1567 -254 1575 -245
rect 1577 -254 1588 -241
rect 1567 -263 1572 -254
rect 1579 -262 1588 -254
rect 1549 -264 1556 -263
rect 1542 -266 1556 -264
rect 1579 -264 1582 -262
rect 1584 -264 1588 -262
rect 1579 -266 1588 -264
rect 1590 -243 1597 -241
rect 1590 -245 1593 -243
rect 1595 -245 1597 -243
rect 1621 -245 1629 -238
rect 1590 -250 1597 -245
rect 1590 -252 1593 -250
rect 1595 -252 1597 -250
rect 1590 -254 1597 -252
rect 1604 -253 1609 -245
rect 1590 -266 1595 -254
rect 1602 -255 1609 -253
rect 1602 -257 1604 -255
rect 1606 -257 1609 -255
rect 1602 -259 1609 -257
rect 1604 -266 1609 -259
rect 1611 -266 1616 -245
rect 1618 -256 1629 -245
rect 1631 -243 1636 -238
rect 1631 -245 1638 -243
rect 1631 -247 1634 -245
rect 1636 -247 1638 -245
rect 1671 -246 1677 -239
rect 1631 -252 1638 -247
rect 1631 -254 1634 -252
rect 1636 -254 1638 -252
rect 1631 -256 1638 -254
rect 1650 -255 1657 -246
rect 1618 -262 1627 -256
rect 1650 -257 1652 -255
rect 1654 -257 1657 -255
rect 1650 -259 1657 -257
rect 1659 -248 1667 -246
rect 1659 -250 1662 -248
rect 1664 -250 1667 -248
rect 1659 -255 1667 -250
rect 1659 -257 1662 -255
rect 1664 -257 1667 -255
rect 1659 -259 1667 -257
rect 1669 -253 1677 -246
rect 1669 -255 1672 -253
rect 1674 -255 1677 -253
rect 1669 -257 1677 -255
rect 1679 -241 1686 -239
rect 1715 -241 1720 -238
rect 1679 -243 1682 -241
rect 1684 -243 1686 -241
rect 1679 -248 1686 -243
rect 1679 -250 1682 -248
rect 1684 -250 1686 -248
rect 1679 -252 1686 -250
rect 1690 -243 1697 -241
rect 1690 -245 1692 -243
rect 1694 -245 1697 -243
rect 1690 -250 1697 -245
rect 1690 -252 1692 -250
rect 1694 -252 1697 -250
rect 1679 -257 1684 -252
rect 1690 -254 1697 -252
rect 1669 -259 1675 -257
rect 1618 -264 1623 -262
rect 1625 -264 1627 -262
rect 1618 -266 1627 -264
rect 1692 -266 1697 -254
rect 1699 -254 1710 -241
rect 1712 -243 1720 -241
rect 1712 -245 1715 -243
rect 1717 -245 1720 -243
rect 1712 -254 1720 -245
rect 1699 -262 1708 -254
rect 1699 -264 1703 -262
rect 1705 -264 1708 -262
rect 1715 -263 1720 -254
rect 1722 -263 1727 -238
rect 1729 -255 1745 -238
rect 1729 -257 1738 -255
rect 1740 -257 1745 -255
rect 1729 -262 1745 -257
rect 1729 -263 1738 -262
rect 1699 -266 1708 -264
rect 1731 -264 1738 -263
rect 1740 -264 1745 -262
rect 1731 -266 1745 -264
rect 1747 -247 1755 -238
rect 1747 -249 1750 -247
rect 1752 -249 1755 -247
rect 1747 -254 1755 -249
rect 1747 -256 1750 -254
rect 1752 -256 1755 -254
rect 1747 -266 1755 -256
rect 1757 -255 1765 -238
rect 1757 -257 1760 -255
rect 1762 -257 1765 -255
rect 1757 -262 1765 -257
rect 1757 -264 1760 -262
rect 1762 -264 1765 -262
rect 1757 -266 1765 -264
rect 1767 -240 1774 -238
rect 1767 -242 1770 -240
rect 1772 -242 1774 -240
rect 1767 -247 1774 -242
rect 1767 -249 1770 -247
rect 1772 -249 1774 -247
rect 1767 -251 1774 -249
rect 1780 -240 1787 -238
rect 1780 -242 1782 -240
rect 1784 -242 1787 -240
rect 1780 -247 1787 -242
rect 1780 -249 1782 -247
rect 1784 -249 1787 -247
rect 1780 -251 1787 -249
rect 1767 -266 1772 -251
rect 1782 -266 1787 -251
rect 1789 -255 1797 -238
rect 1789 -257 1792 -255
rect 1794 -257 1797 -255
rect 1789 -262 1797 -257
rect 1789 -264 1792 -262
rect 1794 -264 1797 -262
rect 1789 -266 1797 -264
rect 1799 -247 1807 -238
rect 1799 -249 1802 -247
rect 1804 -249 1807 -247
rect 1799 -254 1807 -249
rect 1799 -256 1802 -254
rect 1804 -256 1807 -254
rect 1799 -266 1807 -256
rect 1809 -255 1825 -238
rect 1809 -257 1814 -255
rect 1816 -257 1825 -255
rect 1809 -262 1825 -257
rect 1809 -264 1814 -262
rect 1816 -263 1825 -262
rect 1827 -263 1832 -238
rect 1834 -241 1839 -238
rect 1834 -243 1842 -241
rect 1834 -245 1837 -243
rect 1839 -245 1842 -243
rect 1834 -254 1842 -245
rect 1844 -254 1855 -241
rect 1834 -263 1839 -254
rect 1846 -262 1855 -254
rect 1816 -264 1823 -263
rect 1809 -266 1823 -264
rect 1846 -264 1849 -262
rect 1851 -264 1855 -262
rect 1846 -266 1855 -264
rect 1857 -243 1864 -241
rect 1857 -245 1860 -243
rect 1862 -245 1864 -243
rect 1888 -245 1896 -238
rect 1857 -250 1864 -245
rect 1857 -252 1860 -250
rect 1862 -252 1864 -250
rect 1857 -254 1864 -252
rect 1871 -253 1876 -245
rect 1857 -266 1862 -254
rect 1869 -255 1876 -253
rect 1869 -257 1871 -255
rect 1873 -257 1876 -255
rect 1869 -259 1876 -257
rect 1871 -266 1876 -259
rect 1878 -266 1883 -245
rect 1885 -256 1896 -245
rect 1898 -243 1903 -238
rect 1920 -241 1927 -239
rect 1920 -243 1922 -241
rect 1924 -243 1927 -241
rect 1898 -245 1905 -243
rect 1920 -245 1927 -243
rect 1898 -247 1901 -245
rect 1903 -247 1905 -245
rect 1898 -252 1905 -247
rect 1898 -254 1901 -252
rect 1903 -254 1905 -252
rect 1898 -256 1905 -254
rect 1885 -262 1894 -256
rect 1885 -264 1890 -262
rect 1892 -264 1894 -262
rect 1885 -266 1894 -264
rect 1922 -266 1927 -245
rect 1929 -255 1943 -239
rect 1929 -257 1932 -255
rect 1934 -257 1943 -255
rect 1945 -241 1953 -239
rect 1945 -243 1948 -241
rect 1950 -243 1953 -241
rect 1945 -248 1953 -243
rect 1945 -250 1948 -248
rect 1950 -250 1953 -248
rect 1945 -257 1953 -250
rect 1955 -248 1963 -239
rect 1955 -250 1958 -248
rect 1960 -250 1963 -248
rect 1955 -257 1963 -250
rect 1929 -262 1941 -257
rect 1929 -264 1932 -262
rect 1934 -264 1941 -262
rect 1929 -266 1941 -264
rect 1958 -266 1963 -257
rect 1965 -254 1970 -239
rect 2001 -241 2006 -238
rect 1976 -243 1983 -241
rect 1976 -245 1978 -243
rect 1980 -245 1983 -243
rect 1976 -250 1983 -245
rect 1976 -252 1978 -250
rect 1980 -252 1983 -250
rect 1976 -254 1983 -252
rect 1965 -256 1972 -254
rect 1965 -258 1968 -256
rect 1970 -258 1972 -256
rect 1965 -260 1972 -258
rect 1965 -266 1970 -260
rect 1978 -266 1983 -254
rect 1985 -254 1996 -241
rect 1998 -243 2006 -241
rect 1998 -245 2001 -243
rect 2003 -245 2006 -243
rect 1998 -254 2006 -245
rect 1985 -262 1994 -254
rect 1985 -264 1989 -262
rect 1991 -264 1994 -262
rect 2001 -263 2006 -254
rect 2008 -263 2013 -238
rect 2015 -255 2031 -238
rect 2015 -257 2024 -255
rect 2026 -257 2031 -255
rect 2015 -262 2031 -257
rect 2015 -263 2024 -262
rect 1985 -266 1994 -264
rect 2017 -264 2024 -263
rect 2026 -264 2031 -262
rect 2017 -266 2031 -264
rect 2033 -247 2041 -238
rect 2033 -249 2036 -247
rect 2038 -249 2041 -247
rect 2033 -254 2041 -249
rect 2033 -256 2036 -254
rect 2038 -256 2041 -254
rect 2033 -266 2041 -256
rect 2043 -255 2051 -238
rect 2043 -257 2046 -255
rect 2048 -257 2051 -255
rect 2043 -262 2051 -257
rect 2043 -264 2046 -262
rect 2048 -264 2051 -262
rect 2043 -266 2051 -264
rect 2053 -240 2060 -238
rect 2053 -242 2056 -240
rect 2058 -242 2060 -240
rect 2053 -247 2060 -242
rect 2053 -249 2056 -247
rect 2058 -249 2060 -247
rect 2053 -251 2060 -249
rect 2066 -240 2073 -238
rect 2066 -242 2068 -240
rect 2070 -242 2073 -240
rect 2066 -247 2073 -242
rect 2066 -249 2068 -247
rect 2070 -249 2073 -247
rect 2066 -251 2073 -249
rect 2053 -266 2058 -251
rect 2068 -266 2073 -251
rect 2075 -255 2083 -238
rect 2075 -257 2078 -255
rect 2080 -257 2083 -255
rect 2075 -262 2083 -257
rect 2075 -264 2078 -262
rect 2080 -264 2083 -262
rect 2075 -266 2083 -264
rect 2085 -247 2093 -238
rect 2085 -249 2088 -247
rect 2090 -249 2093 -247
rect 2085 -254 2093 -249
rect 2085 -256 2088 -254
rect 2090 -256 2093 -254
rect 2085 -266 2093 -256
rect 2095 -255 2111 -238
rect 2095 -257 2100 -255
rect 2102 -257 2111 -255
rect 2095 -262 2111 -257
rect 2095 -264 2100 -262
rect 2102 -263 2111 -262
rect 2113 -263 2118 -238
rect 2120 -241 2125 -238
rect 2120 -243 2128 -241
rect 2120 -245 2123 -243
rect 2125 -245 2128 -243
rect 2120 -254 2128 -245
rect 2130 -254 2141 -241
rect 2120 -263 2125 -254
rect 2132 -262 2141 -254
rect 2102 -264 2109 -263
rect 2095 -266 2109 -264
rect 2132 -264 2135 -262
rect 2137 -264 2141 -262
rect 2132 -266 2141 -264
rect 2143 -243 2150 -241
rect 2143 -245 2146 -243
rect 2148 -245 2150 -243
rect 2174 -245 2182 -238
rect 2143 -250 2150 -245
rect 2143 -252 2146 -250
rect 2148 -252 2150 -250
rect 2143 -254 2150 -252
rect 2157 -253 2162 -245
rect 2143 -266 2148 -254
rect 2155 -255 2162 -253
rect 2155 -257 2157 -255
rect 2159 -257 2162 -255
rect 2155 -259 2162 -257
rect 2157 -266 2162 -259
rect 2164 -266 2169 -245
rect 2171 -256 2182 -245
rect 2184 -243 2189 -238
rect 2199 -240 2206 -238
rect 2199 -242 2201 -240
rect 2203 -242 2206 -240
rect 2184 -245 2191 -243
rect 2199 -244 2206 -242
rect 2184 -247 2187 -245
rect 2189 -247 2191 -245
rect 2201 -246 2206 -244
rect 2208 -246 2214 -238
rect 2184 -252 2191 -247
rect 2184 -254 2187 -252
rect 2189 -254 2191 -252
rect 2184 -256 2191 -254
rect 2210 -250 2214 -246
rect 2267 -240 2274 -238
rect 2267 -242 2269 -240
rect 2271 -242 2274 -240
rect 2267 -244 2274 -242
rect 2269 -246 2274 -244
rect 2276 -246 2282 -238
rect 2245 -250 2250 -248
rect 2210 -254 2216 -250
rect 2171 -262 2180 -256
rect 2171 -264 2176 -262
rect 2178 -264 2180 -262
rect 2209 -262 2216 -254
rect 2171 -266 2180 -264
rect 2209 -264 2211 -262
rect 2213 -264 2216 -262
rect 2209 -266 2216 -264
rect 2218 -266 2223 -250
rect 2225 -252 2233 -250
rect 2225 -254 2228 -252
rect 2230 -254 2233 -252
rect 2225 -266 2233 -254
rect 2235 -266 2240 -250
rect 2242 -262 2250 -250
rect 2242 -264 2245 -262
rect 2247 -264 2250 -262
rect 2242 -266 2250 -264
rect 2252 -253 2257 -248
rect 2278 -250 2282 -246
rect 2313 -250 2318 -248
rect 2252 -255 2259 -253
rect 2278 -254 2284 -250
rect 2252 -257 2255 -255
rect 2257 -257 2259 -255
rect 2252 -259 2259 -257
rect 2252 -266 2257 -259
rect 2277 -262 2284 -254
rect 2277 -264 2279 -262
rect 2281 -264 2284 -262
rect 2277 -266 2284 -264
rect 2286 -266 2291 -250
rect 2293 -252 2301 -250
rect 2293 -254 2296 -252
rect 2298 -254 2301 -252
rect 2293 -266 2301 -254
rect 2303 -266 2308 -250
rect 2310 -262 2318 -250
rect 2310 -264 2313 -262
rect 2315 -264 2318 -262
rect 2310 -266 2318 -264
rect 2320 -253 2325 -248
rect 2320 -255 2327 -253
rect 2320 -257 2323 -255
rect 2325 -257 2327 -255
rect 2320 -259 2327 -257
rect 2320 -266 2325 -259
<< alu1 >>
rect 4 303 2331 304
rect 4 301 2320 303
rect 2322 301 2331 303
rect 4 299 2331 301
rect 4 297 39 299
rect 41 297 79 299
rect 81 297 298 299
rect 300 297 346 299
rect 348 297 565 299
rect 567 297 613 299
rect 615 297 832 299
rect 834 297 880 299
rect 882 297 1099 299
rect 1101 297 1147 299
rect 1149 297 1366 299
rect 1368 297 1414 299
rect 1416 297 1633 299
rect 1635 297 1681 299
rect 1683 297 1900 299
rect 1902 297 1948 299
rect 1950 297 2186 299
rect 2188 297 2331 299
rect 4 296 2331 297
rect 8 276 12 283
rect 39 282 44 284
rect 8 274 9 276
rect 11 274 12 276
rect 8 273 21 274
rect 8 271 13 273
rect 15 271 21 273
rect 8 270 21 271
rect 15 265 29 266
rect 15 263 23 265
rect 25 263 29 265
rect 15 262 29 263
rect 39 280 40 282
rect 42 280 44 282
rect 39 275 44 280
rect 39 273 40 275
rect 42 273 44 275
rect 39 271 44 273
rect 15 253 20 262
rect 40 270 44 271
rect 48 274 52 283
rect 299 290 303 291
rect 290 286 303 290
rect 88 284 93 286
rect 79 282 84 284
rect 48 273 61 274
rect 48 271 53 273
rect 55 271 61 273
rect 48 270 61 271
rect 40 268 41 270
rect 43 268 44 270
rect 40 251 44 268
rect 55 265 69 266
rect 55 263 63 265
rect 65 263 69 265
rect 55 262 69 263
rect 79 280 80 282
rect 82 280 84 282
rect 79 275 84 280
rect 79 273 80 275
rect 82 273 84 275
rect 79 271 84 273
rect 55 259 60 262
rect 55 257 57 259
rect 59 257 60 259
rect 55 253 60 257
rect 80 265 84 271
rect 80 263 81 265
rect 83 263 84 265
rect 32 249 40 251
rect 42 249 44 251
rect 80 251 84 263
rect 32 245 44 249
rect 72 249 80 251
rect 82 249 84 251
rect 72 245 84 249
rect 88 282 90 284
rect 92 282 93 284
rect 88 277 93 282
rect 88 275 90 277
rect 92 275 93 277
rect 88 273 93 275
rect 88 257 92 273
rect 119 273 157 274
rect 119 271 121 273
rect 123 271 157 273
rect 119 270 157 271
rect 119 267 124 270
rect 116 265 124 267
rect 116 263 117 265
rect 119 263 124 265
rect 116 261 124 263
rect 134 265 149 266
rect 134 263 136 265
rect 138 263 139 265
rect 141 263 143 265
rect 145 263 149 265
rect 134 262 149 263
rect 88 255 89 257
rect 91 255 92 257
rect 88 251 92 255
rect 88 249 93 251
rect 136 253 140 262
rect 167 281 173 283
rect 167 279 168 281
rect 170 279 173 281
rect 167 274 173 279
rect 167 272 168 274
rect 170 272 173 274
rect 167 270 173 272
rect 169 265 173 270
rect 169 263 170 265
rect 172 263 173 265
rect 169 250 173 263
rect 88 247 90 249
rect 92 247 93 249
rect 88 245 93 247
rect 167 249 173 250
rect 167 247 168 249
rect 170 247 173 249
rect 167 246 173 247
rect 177 281 183 283
rect 257 284 262 286
rect 257 282 258 284
rect 260 282 262 284
rect 177 279 180 281
rect 182 279 183 281
rect 177 278 183 279
rect 177 276 180 278
rect 182 276 183 278
rect 177 274 183 276
rect 177 272 180 274
rect 182 272 183 274
rect 177 270 183 272
rect 177 250 181 270
rect 193 273 231 274
rect 193 271 210 273
rect 212 271 231 273
rect 193 270 231 271
rect 226 267 231 270
rect 201 265 216 266
rect 201 263 205 265
rect 207 263 212 265
rect 214 263 216 265
rect 201 262 216 263
rect 226 265 234 267
rect 226 263 231 265
rect 233 263 234 265
rect 210 257 214 262
rect 226 261 234 263
rect 257 277 262 282
rect 257 275 258 277
rect 260 275 262 277
rect 257 273 262 275
rect 258 271 259 273
rect 261 271 262 273
rect 210 255 211 257
rect 213 255 214 257
rect 210 253 214 255
rect 177 249 183 250
rect 177 247 180 249
rect 182 247 183 249
rect 177 246 183 247
rect 258 251 262 271
rect 267 282 271 283
rect 267 280 268 282
rect 270 280 271 282
rect 267 274 271 280
rect 267 272 288 274
rect 267 270 272 272
rect 274 270 288 272
rect 267 265 288 266
rect 267 263 268 265
rect 270 263 282 265
rect 284 263 288 265
rect 267 262 288 263
rect 301 284 303 286
rect 299 279 303 284
rect 301 277 303 279
rect 267 253 271 262
rect 299 261 303 277
rect 315 274 319 283
rect 566 290 570 291
rect 557 286 570 290
rect 355 284 360 286
rect 346 282 351 284
rect 315 273 328 274
rect 315 271 320 273
rect 322 271 328 273
rect 315 270 328 271
rect 299 259 300 261
rect 302 259 303 261
rect 299 258 303 259
rect 298 256 303 258
rect 298 254 299 256
rect 301 254 303 256
rect 298 252 303 254
rect 322 265 336 266
rect 322 263 330 265
rect 332 263 336 265
rect 322 262 336 263
rect 346 280 347 282
rect 349 280 351 282
rect 346 275 351 280
rect 346 273 347 275
rect 349 273 351 275
rect 346 271 351 273
rect 322 259 327 262
rect 322 257 324 259
rect 326 257 327 259
rect 322 253 327 257
rect 347 265 351 271
rect 347 263 348 265
rect 350 263 351 265
rect 257 249 262 251
rect 347 251 351 263
rect 257 247 258 249
rect 260 247 262 249
rect 257 245 262 247
rect 339 249 347 251
rect 349 249 351 251
rect 339 245 351 249
rect 355 282 357 284
rect 359 282 360 284
rect 355 277 360 282
rect 355 275 357 277
rect 359 275 360 277
rect 355 273 360 275
rect 355 257 359 273
rect 386 273 424 274
rect 386 271 388 273
rect 390 271 424 273
rect 386 270 424 271
rect 386 267 391 270
rect 383 265 391 267
rect 383 263 384 265
rect 386 263 391 265
rect 383 261 391 263
rect 401 265 416 266
rect 401 263 403 265
rect 405 263 406 265
rect 408 263 410 265
rect 412 263 416 265
rect 401 262 416 263
rect 355 255 356 257
rect 358 255 359 257
rect 355 251 359 255
rect 355 249 360 251
rect 403 253 407 262
rect 434 281 440 283
rect 434 279 435 281
rect 437 279 440 281
rect 434 274 440 279
rect 434 272 435 274
rect 437 272 440 274
rect 434 270 440 272
rect 436 265 440 270
rect 436 263 437 265
rect 439 263 440 265
rect 436 250 440 263
rect 355 247 357 249
rect 359 247 360 249
rect 355 245 360 247
rect 434 249 440 250
rect 434 247 435 249
rect 437 247 440 249
rect 434 246 440 247
rect 444 281 450 283
rect 524 284 529 286
rect 524 282 525 284
rect 527 282 529 284
rect 444 279 447 281
rect 449 279 450 281
rect 444 278 450 279
rect 444 276 447 278
rect 449 276 450 278
rect 444 274 450 276
rect 444 272 447 274
rect 449 272 450 274
rect 444 270 450 272
rect 444 250 448 270
rect 460 273 498 274
rect 460 271 477 273
rect 479 271 498 273
rect 460 270 498 271
rect 493 267 498 270
rect 468 265 483 266
rect 468 263 472 265
rect 474 263 479 265
rect 481 263 483 265
rect 468 262 483 263
rect 493 265 501 267
rect 493 263 498 265
rect 500 263 501 265
rect 477 257 481 262
rect 493 261 501 263
rect 524 277 529 282
rect 524 275 525 277
rect 527 275 529 277
rect 524 273 529 275
rect 525 271 526 273
rect 528 271 529 273
rect 477 255 478 257
rect 480 255 481 257
rect 477 253 481 255
rect 444 249 450 250
rect 444 247 447 249
rect 449 247 450 249
rect 444 246 450 247
rect 525 251 529 271
rect 534 282 538 283
rect 534 280 535 282
rect 537 280 538 282
rect 534 274 538 280
rect 534 272 555 274
rect 534 270 539 272
rect 541 270 555 272
rect 534 265 555 266
rect 534 263 535 265
rect 537 263 549 265
rect 551 263 555 265
rect 534 262 555 263
rect 568 284 570 286
rect 566 279 570 284
rect 568 277 570 279
rect 534 253 538 262
rect 566 261 570 277
rect 582 274 586 283
rect 833 290 837 291
rect 824 286 837 290
rect 622 284 627 286
rect 613 282 618 284
rect 582 273 595 274
rect 582 271 587 273
rect 589 271 595 273
rect 582 270 595 271
rect 566 259 567 261
rect 569 259 570 261
rect 566 258 570 259
rect 565 256 570 258
rect 565 254 566 256
rect 568 254 570 256
rect 565 252 570 254
rect 589 265 603 266
rect 589 263 597 265
rect 599 263 603 265
rect 589 262 603 263
rect 613 280 614 282
rect 616 280 618 282
rect 613 275 618 280
rect 613 273 614 275
rect 616 273 618 275
rect 613 271 618 273
rect 589 259 594 262
rect 589 257 591 259
rect 593 257 594 259
rect 589 253 594 257
rect 614 265 618 271
rect 614 263 615 265
rect 617 263 618 265
rect 524 249 529 251
rect 614 251 618 263
rect 524 247 525 249
rect 527 247 529 249
rect 524 245 529 247
rect 606 249 614 251
rect 616 249 618 251
rect 606 245 618 249
rect 622 282 624 284
rect 626 282 627 284
rect 622 277 627 282
rect 622 275 624 277
rect 626 275 627 277
rect 622 273 627 275
rect 622 257 626 273
rect 653 273 691 274
rect 653 271 655 273
rect 657 271 691 273
rect 653 270 691 271
rect 653 267 658 270
rect 650 265 658 267
rect 650 263 651 265
rect 653 263 658 265
rect 650 261 658 263
rect 668 265 683 266
rect 668 263 670 265
rect 672 263 673 265
rect 675 263 677 265
rect 679 263 683 265
rect 668 262 683 263
rect 622 255 623 257
rect 625 255 626 257
rect 622 251 626 255
rect 622 249 627 251
rect 670 253 674 262
rect 701 281 707 283
rect 701 279 702 281
rect 704 279 707 281
rect 701 274 707 279
rect 701 272 702 274
rect 704 272 707 274
rect 701 270 707 272
rect 703 265 707 270
rect 703 263 704 265
rect 706 263 707 265
rect 703 250 707 263
rect 622 247 624 249
rect 626 247 627 249
rect 622 245 627 247
rect 701 249 707 250
rect 701 247 702 249
rect 704 247 707 249
rect 701 246 707 247
rect 711 281 717 283
rect 791 284 796 286
rect 791 282 792 284
rect 794 282 796 284
rect 711 279 714 281
rect 716 279 717 281
rect 711 278 717 279
rect 711 276 714 278
rect 716 276 717 278
rect 711 274 717 276
rect 711 272 714 274
rect 716 272 717 274
rect 711 270 717 272
rect 711 250 715 270
rect 727 273 765 274
rect 727 271 744 273
rect 746 271 765 273
rect 727 270 765 271
rect 760 267 765 270
rect 735 265 750 266
rect 735 263 739 265
rect 741 263 746 265
rect 748 263 750 265
rect 735 262 750 263
rect 760 265 768 267
rect 760 263 765 265
rect 767 263 768 265
rect 744 257 748 262
rect 760 261 768 263
rect 791 277 796 282
rect 791 275 792 277
rect 794 275 796 277
rect 791 273 796 275
rect 744 255 745 257
rect 747 255 748 257
rect 744 253 748 255
rect 711 249 717 250
rect 711 247 714 249
rect 716 247 717 249
rect 711 246 717 247
rect 792 257 796 273
rect 801 282 805 283
rect 801 280 802 282
rect 804 280 805 282
rect 801 274 805 280
rect 801 272 822 274
rect 801 270 806 272
rect 808 270 822 272
rect 792 255 793 257
rect 795 255 796 257
rect 792 251 796 255
rect 801 265 822 266
rect 801 263 802 265
rect 804 263 816 265
rect 818 263 822 265
rect 801 262 822 263
rect 835 284 837 286
rect 833 279 837 284
rect 835 277 837 279
rect 801 253 805 262
rect 833 261 837 277
rect 849 274 853 283
rect 1100 290 1104 291
rect 1091 286 1104 290
rect 889 284 894 286
rect 880 282 885 284
rect 849 273 862 274
rect 849 271 854 273
rect 856 271 862 273
rect 849 270 862 271
rect 833 259 834 261
rect 836 259 837 261
rect 833 258 837 259
rect 832 256 837 258
rect 832 254 833 256
rect 835 254 837 256
rect 832 252 837 254
rect 856 265 870 266
rect 856 263 864 265
rect 866 263 870 265
rect 856 262 870 263
rect 880 280 881 282
rect 883 280 885 282
rect 880 275 885 280
rect 880 273 881 275
rect 883 273 885 275
rect 880 271 885 273
rect 856 259 861 262
rect 856 257 858 259
rect 860 257 861 259
rect 856 253 861 257
rect 881 265 885 271
rect 881 263 882 265
rect 884 263 885 265
rect 791 249 796 251
rect 881 251 885 263
rect 791 247 792 249
rect 794 247 796 249
rect 791 245 796 247
rect 873 249 881 251
rect 883 249 885 251
rect 873 245 885 249
rect 889 282 891 284
rect 893 282 894 284
rect 889 277 894 282
rect 889 275 891 277
rect 893 275 894 277
rect 889 273 894 275
rect 889 257 893 273
rect 920 273 958 274
rect 920 271 922 273
rect 924 271 958 273
rect 920 270 958 271
rect 920 267 925 270
rect 917 265 925 267
rect 917 263 918 265
rect 920 263 925 265
rect 917 261 925 263
rect 935 265 950 266
rect 935 263 937 265
rect 939 263 940 265
rect 942 263 944 265
rect 946 263 950 265
rect 935 262 950 263
rect 889 255 890 257
rect 892 255 893 257
rect 889 251 893 255
rect 889 249 894 251
rect 937 253 941 262
rect 968 281 974 283
rect 968 279 969 281
rect 971 279 974 281
rect 968 274 974 279
rect 968 272 969 274
rect 971 272 974 274
rect 968 270 974 272
rect 970 265 974 270
rect 970 263 971 265
rect 973 263 974 265
rect 970 250 974 263
rect 889 247 891 249
rect 893 247 894 249
rect 889 245 894 247
rect 968 249 974 250
rect 968 247 969 249
rect 971 247 974 249
rect 968 246 974 247
rect 978 281 984 283
rect 1058 284 1063 286
rect 1058 282 1059 284
rect 1061 282 1063 284
rect 978 279 981 281
rect 983 279 984 281
rect 978 278 984 279
rect 978 276 981 278
rect 983 276 984 278
rect 978 274 984 276
rect 978 272 981 274
rect 983 272 984 274
rect 978 270 984 272
rect 978 250 982 270
rect 994 273 1032 274
rect 994 271 1011 273
rect 1013 271 1032 273
rect 994 270 1032 271
rect 1027 267 1032 270
rect 1002 265 1017 266
rect 1002 263 1006 265
rect 1008 263 1013 265
rect 1015 263 1017 265
rect 1002 262 1017 263
rect 1027 265 1035 267
rect 1027 263 1032 265
rect 1034 263 1035 265
rect 1011 257 1015 262
rect 1027 261 1035 263
rect 1058 277 1063 282
rect 1058 275 1059 277
rect 1061 275 1063 277
rect 1058 273 1063 275
rect 1011 255 1012 257
rect 1014 255 1015 257
rect 1011 253 1015 255
rect 978 249 984 250
rect 978 247 981 249
rect 983 247 984 249
rect 978 246 984 247
rect 1059 257 1063 273
rect 1068 282 1072 283
rect 1068 280 1069 282
rect 1071 280 1072 282
rect 1068 274 1072 280
rect 1068 272 1089 274
rect 1068 270 1073 272
rect 1075 270 1089 272
rect 1059 255 1060 257
rect 1062 255 1063 257
rect 1059 251 1063 255
rect 1068 265 1089 266
rect 1068 263 1069 265
rect 1071 263 1083 265
rect 1085 263 1089 265
rect 1068 262 1089 263
rect 1102 284 1104 286
rect 1100 279 1104 284
rect 1102 277 1104 279
rect 1068 253 1072 262
rect 1100 261 1104 277
rect 1116 274 1120 283
rect 1367 290 1371 291
rect 1358 286 1371 290
rect 1156 284 1161 286
rect 1147 282 1152 284
rect 1116 273 1129 274
rect 1116 271 1121 273
rect 1123 271 1129 273
rect 1116 270 1129 271
rect 1100 259 1101 261
rect 1103 259 1104 261
rect 1100 258 1104 259
rect 1099 256 1104 258
rect 1099 254 1100 256
rect 1102 254 1104 256
rect 1099 252 1104 254
rect 1123 265 1137 266
rect 1123 263 1131 265
rect 1133 263 1137 265
rect 1123 262 1137 263
rect 1147 280 1148 282
rect 1150 280 1152 282
rect 1147 275 1152 280
rect 1147 273 1148 275
rect 1150 273 1152 275
rect 1147 271 1152 273
rect 1123 259 1128 262
rect 1123 257 1125 259
rect 1127 257 1128 259
rect 1123 253 1128 257
rect 1148 265 1152 271
rect 1148 263 1149 265
rect 1151 263 1152 265
rect 1058 249 1063 251
rect 1148 251 1152 263
rect 1058 247 1059 249
rect 1061 247 1063 249
rect 1058 245 1063 247
rect 1140 249 1148 251
rect 1150 249 1152 251
rect 1140 245 1152 249
rect 1156 282 1158 284
rect 1160 282 1161 284
rect 1156 277 1161 282
rect 1156 275 1158 277
rect 1160 275 1161 277
rect 1156 273 1161 275
rect 1156 257 1160 273
rect 1187 273 1225 274
rect 1187 271 1189 273
rect 1191 271 1225 273
rect 1187 270 1225 271
rect 1187 267 1192 270
rect 1184 265 1192 267
rect 1184 263 1185 265
rect 1187 263 1192 265
rect 1184 261 1192 263
rect 1202 265 1217 266
rect 1202 263 1204 265
rect 1206 263 1207 265
rect 1209 263 1211 265
rect 1213 263 1217 265
rect 1202 262 1217 263
rect 1156 255 1157 257
rect 1159 255 1160 257
rect 1156 251 1160 255
rect 1156 249 1161 251
rect 1204 253 1208 262
rect 1235 281 1241 283
rect 1235 279 1236 281
rect 1238 279 1241 281
rect 1235 274 1241 279
rect 1235 272 1236 274
rect 1238 272 1241 274
rect 1235 270 1241 272
rect 1237 265 1241 270
rect 1237 263 1238 265
rect 1240 263 1241 265
rect 1237 250 1241 263
rect 1156 247 1158 249
rect 1160 247 1161 249
rect 1156 245 1161 247
rect 1235 249 1241 250
rect 1235 247 1236 249
rect 1238 247 1241 249
rect 1235 246 1241 247
rect 1245 281 1251 283
rect 1325 284 1330 286
rect 1325 282 1326 284
rect 1328 282 1330 284
rect 1245 279 1248 281
rect 1250 279 1251 281
rect 1245 278 1251 279
rect 1245 276 1248 278
rect 1250 276 1251 278
rect 1245 274 1251 276
rect 1245 272 1248 274
rect 1250 272 1251 274
rect 1245 270 1251 272
rect 1245 250 1249 270
rect 1261 273 1299 274
rect 1261 271 1278 273
rect 1280 271 1299 273
rect 1261 270 1299 271
rect 1294 267 1299 270
rect 1269 265 1284 266
rect 1269 263 1273 265
rect 1275 263 1280 265
rect 1282 263 1284 265
rect 1269 262 1284 263
rect 1294 265 1302 267
rect 1294 263 1299 265
rect 1301 263 1302 265
rect 1278 257 1282 262
rect 1294 261 1302 263
rect 1325 277 1330 282
rect 1325 275 1326 277
rect 1328 275 1330 277
rect 1325 273 1330 275
rect 1278 255 1279 257
rect 1281 255 1282 257
rect 1278 253 1282 255
rect 1245 249 1251 250
rect 1245 247 1248 249
rect 1250 247 1251 249
rect 1245 246 1251 247
rect 1326 254 1330 273
rect 1335 282 1339 283
rect 1335 280 1336 282
rect 1338 280 1339 282
rect 1335 274 1339 280
rect 1335 272 1356 274
rect 1335 270 1340 272
rect 1342 270 1356 272
rect 1326 252 1327 254
rect 1329 252 1330 254
rect 1335 265 1356 266
rect 1335 263 1336 265
rect 1338 263 1350 265
rect 1352 263 1356 265
rect 1335 262 1356 263
rect 1369 284 1371 286
rect 1367 279 1371 284
rect 1369 277 1371 279
rect 1335 253 1339 262
rect 1367 261 1371 277
rect 1383 274 1387 283
rect 1634 290 1638 291
rect 1625 286 1638 290
rect 1423 284 1428 286
rect 1414 282 1419 284
rect 1383 273 1396 274
rect 1383 271 1388 273
rect 1390 271 1396 273
rect 1383 270 1396 271
rect 1367 259 1368 261
rect 1370 259 1371 261
rect 1367 258 1371 259
rect 1366 256 1371 258
rect 1366 254 1367 256
rect 1369 254 1371 256
rect 1366 252 1371 254
rect 1390 265 1404 266
rect 1390 263 1398 265
rect 1400 263 1404 265
rect 1390 262 1404 263
rect 1414 280 1415 282
rect 1417 280 1419 282
rect 1414 275 1419 280
rect 1414 273 1415 275
rect 1417 273 1419 275
rect 1414 271 1419 273
rect 1390 259 1395 262
rect 1390 257 1392 259
rect 1394 257 1395 259
rect 1390 253 1395 257
rect 1415 265 1419 271
rect 1415 263 1416 265
rect 1418 263 1419 265
rect 1326 251 1330 252
rect 1325 249 1330 251
rect 1415 251 1419 263
rect 1325 247 1326 249
rect 1328 247 1330 249
rect 1325 245 1330 247
rect 1407 249 1415 251
rect 1417 249 1419 251
rect 1407 245 1419 249
rect 1423 282 1425 284
rect 1427 282 1428 284
rect 1423 277 1428 282
rect 1423 275 1425 277
rect 1427 275 1428 277
rect 1423 273 1428 275
rect 1423 257 1427 273
rect 1454 273 1492 274
rect 1454 271 1456 273
rect 1458 271 1492 273
rect 1454 270 1492 271
rect 1454 267 1459 270
rect 1451 265 1459 267
rect 1451 263 1452 265
rect 1454 263 1459 265
rect 1451 261 1459 263
rect 1469 265 1484 266
rect 1469 263 1471 265
rect 1473 263 1474 265
rect 1476 263 1478 265
rect 1480 263 1484 265
rect 1469 262 1484 263
rect 1423 255 1424 257
rect 1426 255 1427 257
rect 1423 251 1427 255
rect 1423 249 1428 251
rect 1471 253 1475 262
rect 1502 281 1508 283
rect 1502 279 1503 281
rect 1505 279 1508 281
rect 1502 274 1508 279
rect 1502 272 1503 274
rect 1505 272 1508 274
rect 1502 270 1508 272
rect 1504 265 1508 270
rect 1504 263 1505 265
rect 1507 263 1508 265
rect 1504 250 1508 263
rect 1423 247 1425 249
rect 1427 247 1428 249
rect 1423 245 1428 247
rect 1502 249 1508 250
rect 1502 247 1503 249
rect 1505 247 1508 249
rect 1502 246 1508 247
rect 1512 281 1518 283
rect 1592 284 1597 286
rect 1592 282 1593 284
rect 1595 282 1597 284
rect 1512 279 1515 281
rect 1517 279 1518 281
rect 1512 278 1518 279
rect 1512 276 1515 278
rect 1517 276 1518 278
rect 1512 274 1518 276
rect 1512 272 1515 274
rect 1517 272 1518 274
rect 1512 270 1518 272
rect 1512 250 1516 270
rect 1528 273 1566 274
rect 1528 271 1545 273
rect 1547 271 1566 273
rect 1528 270 1566 271
rect 1561 267 1566 270
rect 1536 265 1551 266
rect 1536 263 1540 265
rect 1542 263 1547 265
rect 1549 263 1551 265
rect 1536 262 1551 263
rect 1561 265 1569 267
rect 1561 263 1566 265
rect 1568 263 1569 265
rect 1545 257 1549 262
rect 1561 261 1569 263
rect 1592 277 1597 282
rect 1592 275 1593 277
rect 1595 275 1597 277
rect 1592 273 1597 275
rect 1545 255 1546 257
rect 1548 255 1549 257
rect 1545 253 1549 255
rect 1512 249 1518 250
rect 1512 247 1515 249
rect 1517 247 1518 249
rect 1512 246 1518 247
rect 1593 254 1597 273
rect 1602 282 1606 283
rect 1602 280 1603 282
rect 1605 280 1606 282
rect 1602 274 1606 280
rect 1602 272 1623 274
rect 1602 270 1607 272
rect 1609 270 1623 272
rect 1593 252 1594 254
rect 1596 252 1597 254
rect 1602 265 1623 266
rect 1602 263 1603 265
rect 1605 263 1617 265
rect 1619 263 1623 265
rect 1602 262 1623 263
rect 1636 284 1638 286
rect 1634 279 1638 284
rect 1636 277 1638 279
rect 1602 253 1606 262
rect 1634 261 1638 277
rect 1650 274 1654 283
rect 1901 290 1905 291
rect 1892 286 1905 290
rect 1690 284 1695 286
rect 1681 282 1686 284
rect 1650 273 1663 274
rect 1650 271 1655 273
rect 1657 271 1663 273
rect 1650 270 1663 271
rect 1634 259 1635 261
rect 1637 259 1638 261
rect 1634 258 1638 259
rect 1633 256 1638 258
rect 1633 254 1634 256
rect 1636 254 1638 256
rect 1633 252 1638 254
rect 1657 265 1671 266
rect 1657 263 1665 265
rect 1667 263 1671 265
rect 1657 262 1671 263
rect 1681 280 1682 282
rect 1684 280 1686 282
rect 1681 275 1686 280
rect 1681 273 1682 275
rect 1684 273 1686 275
rect 1681 271 1686 273
rect 1657 259 1662 262
rect 1657 257 1659 259
rect 1661 257 1662 259
rect 1657 253 1662 257
rect 1682 265 1686 271
rect 1682 263 1683 265
rect 1685 263 1686 265
rect 1593 251 1597 252
rect 1592 249 1597 251
rect 1682 251 1686 263
rect 1592 247 1593 249
rect 1595 247 1597 249
rect 1592 245 1597 247
rect 1674 249 1682 251
rect 1684 249 1686 251
rect 1674 245 1686 249
rect 1690 282 1692 284
rect 1694 282 1695 284
rect 1690 277 1695 282
rect 1690 275 1692 277
rect 1694 275 1695 277
rect 1690 273 1695 275
rect 1690 257 1694 273
rect 1721 273 1759 274
rect 1721 271 1723 273
rect 1725 271 1759 273
rect 1721 270 1759 271
rect 1721 267 1726 270
rect 1718 265 1726 267
rect 1718 263 1719 265
rect 1721 263 1726 265
rect 1718 261 1726 263
rect 1736 265 1751 266
rect 1736 263 1738 265
rect 1740 263 1741 265
rect 1743 263 1745 265
rect 1747 263 1751 265
rect 1736 262 1751 263
rect 1690 255 1691 257
rect 1693 255 1694 257
rect 1690 251 1694 255
rect 1690 249 1695 251
rect 1738 253 1742 262
rect 1769 281 1775 283
rect 1769 279 1770 281
rect 1772 279 1775 281
rect 1769 274 1775 279
rect 1769 272 1770 274
rect 1772 272 1775 274
rect 1769 270 1775 272
rect 1771 265 1775 270
rect 1771 263 1772 265
rect 1774 263 1775 265
rect 1771 250 1775 263
rect 1690 247 1692 249
rect 1694 247 1695 249
rect 1690 245 1695 247
rect 1769 249 1775 250
rect 1769 247 1770 249
rect 1772 247 1775 249
rect 1769 246 1775 247
rect 1779 281 1785 283
rect 1859 284 1864 286
rect 1859 282 1860 284
rect 1862 282 1864 284
rect 1779 279 1782 281
rect 1784 279 1785 281
rect 1779 278 1785 279
rect 1779 276 1782 278
rect 1784 276 1785 278
rect 1779 274 1785 276
rect 1779 272 1782 274
rect 1784 272 1785 274
rect 1779 270 1785 272
rect 1779 250 1783 270
rect 1795 273 1833 274
rect 1795 271 1812 273
rect 1814 271 1833 273
rect 1795 270 1833 271
rect 1828 267 1833 270
rect 1803 265 1818 266
rect 1803 263 1807 265
rect 1809 263 1814 265
rect 1816 263 1818 265
rect 1803 262 1818 263
rect 1828 265 1836 267
rect 1828 263 1833 265
rect 1835 263 1836 265
rect 1812 257 1816 262
rect 1828 261 1836 263
rect 1859 277 1864 282
rect 1859 275 1860 277
rect 1862 275 1864 277
rect 1859 273 1864 275
rect 1860 271 1861 273
rect 1863 271 1864 273
rect 1812 255 1813 257
rect 1815 255 1816 257
rect 1812 253 1816 255
rect 1779 249 1785 250
rect 1779 247 1782 249
rect 1784 247 1785 249
rect 1779 246 1785 247
rect 1860 251 1864 271
rect 1869 282 1873 283
rect 1869 280 1870 282
rect 1872 280 1873 282
rect 1869 274 1873 280
rect 1869 272 1890 274
rect 1869 270 1874 272
rect 1876 270 1890 272
rect 1869 265 1890 266
rect 1869 263 1870 265
rect 1872 263 1884 265
rect 1886 263 1890 265
rect 1869 262 1890 263
rect 1903 284 1905 286
rect 1901 279 1905 284
rect 1903 277 1905 279
rect 1869 253 1873 262
rect 1901 261 1905 277
rect 1912 285 1924 291
rect 1912 273 1917 285
rect 2187 290 2191 291
rect 2178 286 2191 290
rect 1976 284 1981 286
rect 1912 271 1914 273
rect 1916 271 1917 273
rect 1912 269 1917 271
rect 1901 259 1902 261
rect 1904 259 1905 261
rect 1901 258 1905 259
rect 1900 256 1905 258
rect 1900 254 1901 256
rect 1903 254 1905 256
rect 1900 252 1905 254
rect 1928 260 1933 267
rect 1956 282 1972 283
rect 1956 280 1958 282
rect 1960 280 1972 282
rect 1956 278 1972 280
rect 1968 273 1972 278
rect 1968 271 1969 273
rect 1971 271 1972 273
rect 1928 259 1930 260
rect 1920 258 1930 259
rect 1932 258 1933 260
rect 1920 256 1933 258
rect 1920 254 1925 256
rect 1927 254 1933 256
rect 1920 253 1933 254
rect 1859 249 1864 251
rect 1968 250 1972 271
rect 1859 247 1860 249
rect 1862 247 1864 249
rect 1859 245 1864 247
rect 1948 249 1972 250
rect 1948 247 1950 249
rect 1952 247 1972 249
rect 1948 246 1972 247
rect 1976 282 1978 284
rect 1980 282 1981 284
rect 1976 277 1981 282
rect 1976 275 1978 277
rect 1980 275 1981 277
rect 1976 273 1981 275
rect 1976 257 1980 273
rect 2007 273 2045 274
rect 2007 271 2018 273
rect 2020 271 2045 273
rect 2007 270 2045 271
rect 2007 267 2012 270
rect 2004 265 2012 267
rect 2004 263 2005 265
rect 2007 263 2012 265
rect 2004 261 2012 263
rect 2022 265 2037 266
rect 2022 263 2024 265
rect 2026 263 2031 265
rect 2033 263 2037 265
rect 2022 262 2037 263
rect 1976 255 1977 257
rect 1979 255 1980 257
rect 1976 251 1980 255
rect 1976 249 1981 251
rect 2024 253 2028 262
rect 2055 281 2061 283
rect 2055 279 2056 281
rect 2058 279 2061 281
rect 2055 274 2061 279
rect 2055 272 2056 274
rect 2058 272 2061 274
rect 2055 270 2061 272
rect 2057 265 2061 270
rect 2057 263 2058 265
rect 2060 263 2061 265
rect 2057 250 2061 263
rect 1976 247 1978 249
rect 1980 247 1981 249
rect 1976 245 1981 247
rect 2055 249 2061 250
rect 2055 247 2056 249
rect 2058 247 2061 249
rect 2055 246 2061 247
rect 2065 281 2071 283
rect 2145 284 2150 286
rect 2145 282 2146 284
rect 2148 282 2150 284
rect 2065 279 2068 281
rect 2070 279 2071 281
rect 2065 278 2071 279
rect 2065 276 2068 278
rect 2070 276 2071 278
rect 2065 274 2071 276
rect 2065 272 2068 274
rect 2070 272 2071 274
rect 2065 270 2071 272
rect 2065 250 2069 270
rect 2081 273 2119 274
rect 2081 271 2100 273
rect 2102 271 2119 273
rect 2081 270 2119 271
rect 2114 267 2119 270
rect 2089 265 2104 266
rect 2089 263 2093 265
rect 2095 263 2100 265
rect 2102 263 2104 265
rect 2089 262 2104 263
rect 2114 265 2122 267
rect 2114 263 2119 265
rect 2121 263 2122 265
rect 2098 257 2102 262
rect 2114 261 2122 263
rect 2145 277 2150 282
rect 2145 275 2146 277
rect 2148 275 2150 277
rect 2145 273 2150 275
rect 2098 255 2099 257
rect 2101 255 2102 257
rect 2098 253 2102 255
rect 2065 249 2071 250
rect 2065 247 2068 249
rect 2070 247 2071 249
rect 2065 246 2071 247
rect 2146 257 2150 273
rect 2155 278 2159 283
rect 2155 276 2156 278
rect 2158 276 2159 278
rect 2155 274 2159 276
rect 2155 272 2176 274
rect 2155 270 2160 272
rect 2162 270 2176 272
rect 2146 255 2147 257
rect 2149 255 2150 257
rect 2146 251 2150 255
rect 2155 265 2176 266
rect 2155 263 2156 265
rect 2158 263 2170 265
rect 2172 263 2176 265
rect 2155 262 2176 263
rect 2189 284 2191 286
rect 2187 279 2191 284
rect 2189 277 2191 279
rect 2199 285 2204 291
rect 2246 289 2259 290
rect 2246 287 2255 289
rect 2257 287 2259 289
rect 2199 283 2201 285
rect 2203 283 2204 285
rect 2246 286 2259 287
rect 2199 282 2204 283
rect 2199 278 2212 282
rect 2155 253 2159 262
rect 2187 261 2191 277
rect 2187 259 2188 261
rect 2190 259 2191 261
rect 2187 258 2191 259
rect 2186 256 2191 258
rect 2186 254 2187 256
rect 2189 254 2191 256
rect 2186 252 2191 254
rect 2145 249 2150 251
rect 2145 247 2146 249
rect 2148 247 2150 249
rect 2213 265 2219 267
rect 2213 263 2214 265
rect 2216 263 2219 265
rect 2213 258 2219 263
rect 2206 257 2219 258
rect 2206 255 2208 257
rect 2210 255 2219 257
rect 2231 273 2243 275
rect 2231 271 2236 273
rect 2238 271 2243 273
rect 2231 270 2243 271
rect 2231 269 2241 270
rect 2239 268 2241 269
rect 2239 261 2243 268
rect 2206 254 2219 255
rect 2255 253 2259 286
rect 2267 285 2272 291
rect 2314 289 2327 290
rect 2314 287 2323 289
rect 2325 287 2327 289
rect 2267 283 2269 285
rect 2271 283 2272 285
rect 2314 286 2327 287
rect 2267 282 2272 283
rect 2267 278 2280 282
rect 2254 251 2259 253
rect 2145 245 2150 247
rect 2254 249 2255 251
rect 2257 249 2259 251
rect 2254 247 2259 249
rect 2281 265 2287 267
rect 2281 263 2282 265
rect 2284 263 2287 265
rect 2281 258 2287 263
rect 2274 257 2287 258
rect 2274 255 2276 257
rect 2278 255 2287 257
rect 2299 274 2311 275
rect 2299 272 2300 274
rect 2302 272 2311 274
rect 2299 270 2311 272
rect 2299 269 2309 270
rect 2307 268 2309 269
rect 2307 261 2311 268
rect 2274 254 2287 255
rect 2323 253 2327 286
rect 2322 251 2327 253
rect 2255 245 2259 247
rect 2322 249 2323 251
rect 2325 249 2327 251
rect 2322 247 2327 249
rect 2323 245 2327 247
rect 4 239 2331 240
rect 4 237 29 239
rect 31 237 39 239
rect 41 237 69 239
rect 71 237 79 239
rect 81 237 298 239
rect 300 237 336 239
rect 338 237 346 239
rect 348 237 565 239
rect 567 237 603 239
rect 605 237 613 239
rect 615 237 832 239
rect 834 237 870 239
rect 872 237 880 239
rect 882 237 1099 239
rect 1101 237 1137 239
rect 1139 237 1147 239
rect 1149 237 1366 239
rect 1368 237 1404 239
rect 1406 237 1414 239
rect 1416 237 1633 239
rect 1635 237 1671 239
rect 1673 237 1681 239
rect 1683 237 1900 239
rect 1902 237 1915 239
rect 1917 237 1968 239
rect 1970 237 2186 239
rect 2188 237 2331 239
rect 4 236 2331 237
rect 4 234 216 236
rect 218 234 483 236
rect 485 234 750 236
rect 752 234 1017 236
rect 1019 234 1284 236
rect 1286 234 1551 236
rect 1553 234 1818 236
rect 1820 234 2331 236
rect 4 233 2331 234
rect 4 231 2276 233
rect 2278 231 2331 233
rect 4 229 2331 231
rect 4 227 2311 229
rect 2313 227 2331 229
rect 4 225 29 227
rect 31 225 39 227
rect 41 225 69 227
rect 71 225 79 227
rect 81 225 298 227
rect 300 225 336 227
rect 338 225 346 227
rect 348 225 565 227
rect 567 225 603 227
rect 605 225 613 227
rect 615 225 832 227
rect 834 225 870 227
rect 872 225 880 227
rect 882 225 1099 227
rect 1101 225 1137 227
rect 1139 225 1147 227
rect 1149 225 1366 227
rect 1368 225 1404 227
rect 1406 225 1414 227
rect 1416 225 1633 227
rect 1635 225 1671 227
rect 1673 225 1681 227
rect 1683 225 1900 227
rect 1902 225 1915 227
rect 1917 225 1968 227
rect 1970 225 2186 227
rect 2188 225 2331 227
rect 4 224 2331 225
rect 15 205 20 211
rect 32 215 44 219
rect 32 213 40 215
rect 42 213 44 215
rect 15 203 17 205
rect 19 203 20 205
rect 15 202 20 203
rect 15 201 29 202
rect 15 199 23 201
rect 25 199 29 201
rect 15 198 29 199
rect 8 193 21 194
rect 8 191 13 193
rect 15 191 21 193
rect 8 190 21 191
rect 8 181 12 190
rect 40 193 44 213
rect 55 202 60 211
rect 72 215 84 219
rect 72 213 80 215
rect 82 213 84 215
rect 55 201 69 202
rect 55 199 63 201
rect 65 199 69 201
rect 55 198 69 199
rect 39 191 41 193
rect 43 191 44 193
rect 39 190 44 191
rect 39 188 40 190
rect 42 188 44 190
rect 39 182 44 188
rect 39 180 40 182
rect 42 180 44 182
rect 48 193 61 194
rect 48 191 53 193
rect 55 191 61 193
rect 48 190 61 191
rect 48 185 52 190
rect 80 201 84 213
rect 80 199 81 201
rect 83 199 84 201
rect 80 193 84 199
rect 48 183 49 185
rect 51 183 52 185
rect 48 181 52 183
rect 79 191 84 193
rect 79 189 80 191
rect 82 189 84 191
rect 79 184 84 189
rect 39 178 44 180
rect 79 182 80 184
rect 82 182 84 184
rect 79 180 84 182
rect 88 217 93 219
rect 88 215 90 217
rect 92 215 93 217
rect 88 213 93 215
rect 88 209 92 213
rect 88 207 89 209
rect 91 207 92 209
rect 88 191 92 207
rect 167 217 173 218
rect 167 215 168 217
rect 170 215 173 217
rect 167 214 173 215
rect 88 189 93 191
rect 88 187 90 189
rect 92 187 93 189
rect 88 182 93 187
rect 116 201 124 203
rect 136 202 140 211
rect 116 199 117 201
rect 119 199 124 201
rect 116 197 124 199
rect 134 201 149 202
rect 134 199 136 201
rect 138 199 139 201
rect 141 199 143 201
rect 145 199 149 201
rect 134 198 149 199
rect 119 194 124 197
rect 169 201 173 214
rect 169 199 170 201
rect 172 199 173 201
rect 119 193 157 194
rect 119 191 134 193
rect 136 191 157 193
rect 119 190 157 191
rect 169 194 173 199
rect 167 192 173 194
rect 167 190 168 192
rect 170 190 173 192
rect 167 185 173 190
rect 167 183 168 185
rect 170 183 173 185
rect 88 180 90 182
rect 92 180 93 182
rect 88 178 93 180
rect 167 181 173 183
rect 177 217 183 218
rect 177 215 180 217
rect 182 215 183 217
rect 177 214 183 215
rect 257 218 264 219
rect 257 217 261 218
rect 257 215 258 217
rect 260 216 261 217
rect 263 216 264 218
rect 260 215 264 216
rect 177 194 181 214
rect 210 209 214 211
rect 210 207 211 209
rect 213 207 214 209
rect 177 192 183 194
rect 177 190 180 192
rect 182 190 183 192
rect 177 188 183 190
rect 177 186 180 188
rect 182 186 183 188
rect 177 185 183 186
rect 177 183 180 185
rect 182 183 183 185
rect 177 181 183 183
rect 210 202 214 207
rect 257 213 264 215
rect 201 201 216 202
rect 201 199 205 201
rect 207 199 212 201
rect 214 199 216 201
rect 201 198 216 199
rect 226 201 234 203
rect 226 199 231 201
rect 233 199 234 201
rect 226 197 234 199
rect 226 196 231 197
rect 226 194 228 196
rect 230 194 231 196
rect 193 190 231 194
rect 258 191 262 213
rect 267 207 271 208
rect 267 205 268 207
rect 270 205 271 207
rect 267 202 271 205
rect 267 201 288 202
rect 267 199 282 201
rect 284 199 288 201
rect 267 198 288 199
rect 298 210 303 212
rect 298 208 299 210
rect 301 208 303 210
rect 298 206 303 208
rect 257 189 262 191
rect 257 187 258 189
rect 260 187 262 189
rect 257 182 262 187
rect 257 180 258 182
rect 260 180 262 182
rect 267 192 272 194
rect 274 192 288 194
rect 267 190 288 192
rect 267 188 271 190
rect 267 186 268 188
rect 270 186 271 188
rect 267 181 271 186
rect 257 178 262 180
rect 299 187 303 206
rect 322 202 327 211
rect 339 215 351 219
rect 339 213 347 215
rect 349 213 351 215
rect 322 201 336 202
rect 322 199 330 201
rect 332 199 336 201
rect 322 198 336 199
rect 301 185 303 187
rect 299 180 303 185
rect 315 193 328 194
rect 315 191 320 193
rect 322 191 328 193
rect 315 190 328 191
rect 315 185 319 190
rect 347 201 351 213
rect 347 199 348 201
rect 350 199 351 201
rect 347 193 351 199
rect 315 183 316 185
rect 318 183 319 185
rect 315 181 319 183
rect 346 191 351 193
rect 346 189 347 191
rect 349 189 351 191
rect 346 184 351 189
rect 301 178 303 180
rect 290 177 303 178
rect 290 175 292 177
rect 294 175 303 177
rect 290 174 303 175
rect 299 173 303 174
rect 346 182 347 184
rect 349 182 351 184
rect 346 180 351 182
rect 355 217 360 219
rect 355 215 357 217
rect 359 215 360 217
rect 355 213 360 215
rect 355 209 359 213
rect 355 207 356 209
rect 358 207 359 209
rect 355 191 359 207
rect 434 217 440 218
rect 434 215 435 217
rect 437 215 440 217
rect 434 214 440 215
rect 355 189 360 191
rect 355 187 357 189
rect 359 187 360 189
rect 355 182 360 187
rect 383 201 391 203
rect 403 202 407 211
rect 383 199 384 201
rect 386 199 391 201
rect 383 197 391 199
rect 401 201 416 202
rect 401 199 403 201
rect 405 199 406 201
rect 408 199 410 201
rect 412 199 416 201
rect 401 198 416 199
rect 386 194 391 197
rect 436 201 440 214
rect 436 199 437 201
rect 439 199 440 201
rect 386 193 424 194
rect 386 191 401 193
rect 403 191 424 193
rect 386 190 424 191
rect 436 194 440 199
rect 434 192 440 194
rect 434 190 435 192
rect 437 190 440 192
rect 434 185 440 190
rect 434 183 435 185
rect 437 183 440 185
rect 355 180 357 182
rect 359 180 360 182
rect 355 178 360 180
rect 434 181 440 183
rect 444 217 450 218
rect 444 215 447 217
rect 449 215 450 217
rect 444 214 450 215
rect 524 218 531 219
rect 524 217 528 218
rect 524 215 525 217
rect 527 216 528 217
rect 530 216 531 218
rect 527 215 531 216
rect 444 194 448 214
rect 477 209 481 211
rect 477 207 478 209
rect 480 207 481 209
rect 444 192 450 194
rect 444 190 447 192
rect 449 190 450 192
rect 444 188 450 190
rect 444 186 447 188
rect 449 186 450 188
rect 444 185 450 186
rect 444 183 447 185
rect 449 183 450 185
rect 444 181 450 183
rect 477 202 481 207
rect 524 213 531 215
rect 468 201 483 202
rect 468 199 472 201
rect 474 199 479 201
rect 481 199 483 201
rect 468 198 483 199
rect 493 201 501 203
rect 493 199 498 201
rect 500 199 501 201
rect 493 197 501 199
rect 493 196 498 197
rect 493 194 495 196
rect 497 194 498 196
rect 460 190 498 194
rect 525 191 529 213
rect 534 207 538 208
rect 534 205 535 207
rect 537 205 538 207
rect 534 202 538 205
rect 534 201 555 202
rect 534 199 549 201
rect 551 199 555 201
rect 534 198 555 199
rect 565 210 570 212
rect 565 208 566 210
rect 568 208 570 210
rect 565 206 570 208
rect 524 189 529 191
rect 524 187 525 189
rect 527 187 529 189
rect 524 182 529 187
rect 524 180 525 182
rect 527 180 529 182
rect 534 192 539 194
rect 541 192 555 194
rect 534 190 555 192
rect 534 188 538 190
rect 534 186 535 188
rect 537 186 538 188
rect 534 181 538 186
rect 524 178 529 180
rect 566 187 570 206
rect 589 202 594 211
rect 606 215 618 219
rect 606 213 614 215
rect 616 213 618 215
rect 589 201 603 202
rect 589 199 597 201
rect 599 199 603 201
rect 589 198 603 199
rect 568 185 570 187
rect 566 180 570 185
rect 582 193 595 194
rect 582 191 587 193
rect 589 191 595 193
rect 582 190 595 191
rect 582 185 586 190
rect 614 201 618 213
rect 614 199 615 201
rect 617 199 618 201
rect 614 193 618 199
rect 582 183 583 185
rect 585 183 586 185
rect 582 181 586 183
rect 613 191 618 193
rect 613 189 614 191
rect 616 189 618 191
rect 613 184 618 189
rect 568 178 570 180
rect 557 177 570 178
rect 557 175 559 177
rect 561 175 570 177
rect 557 174 570 175
rect 566 173 570 174
rect 613 182 614 184
rect 616 182 618 184
rect 613 180 618 182
rect 622 217 627 219
rect 622 215 624 217
rect 626 215 627 217
rect 622 213 627 215
rect 622 209 626 213
rect 622 207 623 209
rect 625 207 626 209
rect 622 191 626 207
rect 701 217 707 218
rect 701 215 702 217
rect 704 215 707 217
rect 701 214 707 215
rect 622 189 627 191
rect 622 187 624 189
rect 626 187 627 189
rect 622 182 627 187
rect 650 201 658 203
rect 670 202 674 211
rect 650 199 651 201
rect 653 199 658 201
rect 650 197 658 199
rect 668 201 683 202
rect 668 199 670 201
rect 672 199 673 201
rect 675 199 677 201
rect 679 199 683 201
rect 668 198 683 199
rect 653 194 658 197
rect 703 201 707 214
rect 703 199 704 201
rect 706 199 707 201
rect 653 193 691 194
rect 653 191 668 193
rect 670 191 691 193
rect 653 190 691 191
rect 703 194 707 199
rect 701 192 707 194
rect 701 190 702 192
rect 704 190 707 192
rect 701 185 707 190
rect 701 183 702 185
rect 704 183 707 185
rect 622 180 624 182
rect 626 180 627 182
rect 622 178 627 180
rect 701 181 707 183
rect 711 217 717 218
rect 711 215 714 217
rect 716 215 717 217
rect 711 214 717 215
rect 791 218 798 219
rect 791 217 795 218
rect 791 215 792 217
rect 794 216 795 217
rect 797 216 798 218
rect 794 215 798 216
rect 711 194 715 214
rect 744 209 748 211
rect 744 207 745 209
rect 747 207 748 209
rect 711 192 717 194
rect 711 190 714 192
rect 716 190 717 192
rect 711 188 717 190
rect 711 186 714 188
rect 716 186 717 188
rect 711 185 717 186
rect 711 183 714 185
rect 716 183 717 185
rect 711 181 717 183
rect 744 202 748 207
rect 791 213 798 215
rect 735 201 750 202
rect 735 199 739 201
rect 741 199 746 201
rect 748 199 750 201
rect 735 198 750 199
rect 760 201 768 203
rect 760 199 765 201
rect 767 199 768 201
rect 760 197 768 199
rect 760 196 765 197
rect 760 194 762 196
rect 764 194 765 196
rect 727 190 765 194
rect 792 191 796 213
rect 801 207 805 208
rect 801 205 802 207
rect 804 205 805 207
rect 801 202 805 205
rect 801 201 822 202
rect 801 199 816 201
rect 818 199 822 201
rect 801 198 822 199
rect 832 210 837 212
rect 832 208 833 210
rect 835 208 837 210
rect 832 206 837 208
rect 791 189 796 191
rect 791 187 792 189
rect 794 187 796 189
rect 791 182 796 187
rect 791 180 792 182
rect 794 180 796 182
rect 801 192 806 194
rect 808 192 822 194
rect 801 190 822 192
rect 801 188 805 190
rect 801 186 802 188
rect 804 186 805 188
rect 801 181 805 186
rect 791 178 796 180
rect 833 187 837 206
rect 856 202 861 211
rect 873 215 885 219
rect 873 213 881 215
rect 883 213 885 215
rect 856 201 870 202
rect 856 199 864 201
rect 866 199 870 201
rect 856 198 870 199
rect 835 185 837 187
rect 833 180 837 185
rect 849 193 862 194
rect 849 191 854 193
rect 856 191 862 193
rect 849 190 862 191
rect 849 185 853 190
rect 881 201 885 213
rect 881 199 882 201
rect 884 199 885 201
rect 881 193 885 199
rect 849 183 850 185
rect 852 183 853 185
rect 849 181 853 183
rect 880 191 885 193
rect 880 189 881 191
rect 883 189 885 191
rect 880 184 885 189
rect 835 178 837 180
rect 824 177 837 178
rect 824 175 826 177
rect 828 175 837 177
rect 824 174 837 175
rect 833 173 837 174
rect 880 182 881 184
rect 883 182 885 184
rect 880 180 885 182
rect 889 217 894 219
rect 889 215 891 217
rect 893 215 894 217
rect 889 213 894 215
rect 889 209 893 213
rect 889 207 890 209
rect 892 207 893 209
rect 889 191 893 207
rect 968 217 974 218
rect 968 215 969 217
rect 971 215 974 217
rect 968 214 974 215
rect 889 189 894 191
rect 889 187 891 189
rect 893 187 894 189
rect 889 182 894 187
rect 917 201 925 203
rect 937 202 941 211
rect 917 199 918 201
rect 920 199 925 201
rect 917 197 925 199
rect 935 201 950 202
rect 935 199 937 201
rect 939 199 940 201
rect 942 199 944 201
rect 946 199 950 201
rect 935 198 950 199
rect 920 194 925 197
rect 970 201 974 214
rect 970 199 971 201
rect 973 199 974 201
rect 920 193 958 194
rect 920 191 935 193
rect 937 191 958 193
rect 920 190 958 191
rect 970 194 974 199
rect 968 192 974 194
rect 968 190 969 192
rect 971 190 974 192
rect 968 185 974 190
rect 968 183 969 185
rect 971 183 974 185
rect 889 180 891 182
rect 893 180 894 182
rect 889 178 894 180
rect 968 181 974 183
rect 978 217 984 218
rect 978 215 981 217
rect 983 215 984 217
rect 978 214 984 215
rect 1058 218 1065 219
rect 1058 217 1062 218
rect 1058 215 1059 217
rect 1061 216 1062 217
rect 1064 216 1065 218
rect 1061 215 1065 216
rect 978 194 982 214
rect 1011 209 1015 211
rect 1011 207 1012 209
rect 1014 207 1015 209
rect 978 192 984 194
rect 978 190 981 192
rect 983 190 984 192
rect 978 188 984 190
rect 978 186 981 188
rect 983 186 984 188
rect 978 185 984 186
rect 978 183 981 185
rect 983 183 984 185
rect 978 181 984 183
rect 1011 202 1015 207
rect 1058 213 1065 215
rect 1002 201 1017 202
rect 1002 199 1006 201
rect 1008 199 1013 201
rect 1015 199 1017 201
rect 1002 198 1017 199
rect 1027 201 1035 203
rect 1027 199 1032 201
rect 1034 199 1035 201
rect 1027 197 1035 199
rect 1027 196 1032 197
rect 1027 194 1029 196
rect 1031 194 1032 196
rect 994 190 1032 194
rect 1059 191 1063 213
rect 1068 207 1072 208
rect 1068 205 1069 207
rect 1071 205 1072 207
rect 1068 202 1072 205
rect 1068 201 1089 202
rect 1068 199 1083 201
rect 1085 199 1089 201
rect 1068 198 1089 199
rect 1099 210 1104 212
rect 1099 208 1100 210
rect 1102 208 1104 210
rect 1099 206 1104 208
rect 1058 189 1063 191
rect 1058 187 1059 189
rect 1061 187 1063 189
rect 1058 182 1063 187
rect 1058 180 1059 182
rect 1061 180 1063 182
rect 1068 192 1073 194
rect 1075 192 1089 194
rect 1068 190 1089 192
rect 1068 188 1072 190
rect 1068 186 1069 188
rect 1071 186 1072 188
rect 1068 181 1072 186
rect 1058 178 1063 180
rect 1100 187 1104 206
rect 1123 202 1128 211
rect 1140 215 1152 219
rect 1140 213 1148 215
rect 1150 213 1152 215
rect 1123 201 1137 202
rect 1123 199 1131 201
rect 1133 199 1137 201
rect 1123 198 1137 199
rect 1102 185 1104 187
rect 1100 180 1104 185
rect 1116 193 1129 194
rect 1116 191 1121 193
rect 1123 191 1129 193
rect 1116 190 1129 191
rect 1116 185 1120 190
rect 1148 201 1152 213
rect 1148 199 1149 201
rect 1151 199 1152 201
rect 1148 193 1152 199
rect 1116 183 1117 185
rect 1119 183 1120 185
rect 1116 181 1120 183
rect 1147 191 1152 193
rect 1147 189 1148 191
rect 1150 189 1152 191
rect 1147 184 1152 189
rect 1102 178 1104 180
rect 1091 177 1104 178
rect 1091 175 1093 177
rect 1095 175 1104 177
rect 1091 174 1104 175
rect 1100 173 1104 174
rect 1147 182 1148 184
rect 1150 182 1152 184
rect 1147 180 1152 182
rect 1156 217 1161 219
rect 1156 215 1158 217
rect 1160 215 1161 217
rect 1156 213 1161 215
rect 1156 209 1160 213
rect 1156 207 1157 209
rect 1159 207 1160 209
rect 1156 191 1160 207
rect 1235 217 1241 218
rect 1235 215 1236 217
rect 1238 215 1241 217
rect 1235 214 1241 215
rect 1156 189 1161 191
rect 1156 187 1158 189
rect 1160 187 1161 189
rect 1156 182 1161 187
rect 1184 201 1192 203
rect 1204 202 1208 211
rect 1184 199 1185 201
rect 1187 199 1192 201
rect 1184 197 1192 199
rect 1202 201 1217 202
rect 1202 199 1204 201
rect 1206 199 1207 201
rect 1209 199 1211 201
rect 1213 199 1217 201
rect 1202 198 1217 199
rect 1187 194 1192 197
rect 1237 201 1241 214
rect 1237 199 1238 201
rect 1240 199 1241 201
rect 1187 193 1225 194
rect 1187 191 1202 193
rect 1204 191 1225 193
rect 1187 190 1225 191
rect 1237 194 1241 199
rect 1235 192 1241 194
rect 1235 190 1236 192
rect 1238 190 1241 192
rect 1235 185 1241 190
rect 1235 183 1236 185
rect 1238 183 1241 185
rect 1156 180 1158 182
rect 1160 180 1161 182
rect 1156 178 1161 180
rect 1235 181 1241 183
rect 1245 217 1251 218
rect 1245 215 1248 217
rect 1250 215 1251 217
rect 1245 214 1251 215
rect 1325 218 1332 219
rect 1325 217 1329 218
rect 1325 215 1326 217
rect 1328 216 1329 217
rect 1331 216 1332 218
rect 1328 215 1332 216
rect 1245 194 1249 214
rect 1278 209 1282 211
rect 1278 207 1279 209
rect 1281 207 1282 209
rect 1245 192 1251 194
rect 1245 190 1248 192
rect 1250 190 1251 192
rect 1245 188 1251 190
rect 1245 186 1248 188
rect 1250 186 1251 188
rect 1245 185 1251 186
rect 1245 183 1248 185
rect 1250 183 1251 185
rect 1245 181 1251 183
rect 1278 202 1282 207
rect 1325 213 1332 215
rect 1269 201 1284 202
rect 1269 199 1273 201
rect 1275 199 1280 201
rect 1282 199 1284 201
rect 1269 198 1284 199
rect 1294 201 1302 203
rect 1294 199 1299 201
rect 1301 199 1302 201
rect 1294 197 1302 199
rect 1294 196 1299 197
rect 1294 194 1296 196
rect 1298 194 1299 196
rect 1261 190 1299 194
rect 1326 191 1330 213
rect 1335 207 1339 208
rect 1335 205 1336 207
rect 1338 205 1339 207
rect 1335 202 1339 205
rect 1335 201 1356 202
rect 1335 199 1350 201
rect 1352 199 1356 201
rect 1335 198 1356 199
rect 1366 210 1371 212
rect 1366 208 1367 210
rect 1369 208 1371 210
rect 1366 206 1371 208
rect 1325 189 1330 191
rect 1325 187 1326 189
rect 1328 187 1330 189
rect 1325 182 1330 187
rect 1325 180 1326 182
rect 1328 180 1330 182
rect 1335 192 1340 194
rect 1342 192 1356 194
rect 1335 190 1356 192
rect 1335 188 1339 190
rect 1335 186 1336 188
rect 1338 186 1339 188
rect 1335 181 1339 186
rect 1325 178 1330 180
rect 1367 187 1371 206
rect 1390 202 1395 211
rect 1407 215 1419 219
rect 1407 213 1415 215
rect 1417 213 1419 215
rect 1390 201 1404 202
rect 1390 199 1398 201
rect 1400 199 1404 201
rect 1390 198 1404 199
rect 1369 185 1371 187
rect 1367 180 1371 185
rect 1383 193 1396 194
rect 1383 191 1388 193
rect 1390 191 1396 193
rect 1383 190 1396 191
rect 1383 185 1387 190
rect 1415 201 1419 213
rect 1415 199 1416 201
rect 1418 199 1419 201
rect 1415 193 1419 199
rect 1383 183 1384 185
rect 1386 183 1387 185
rect 1383 181 1387 183
rect 1414 191 1419 193
rect 1414 189 1415 191
rect 1417 189 1419 191
rect 1414 184 1419 189
rect 1369 178 1371 180
rect 1358 177 1371 178
rect 1358 175 1360 177
rect 1362 175 1371 177
rect 1358 174 1371 175
rect 1367 173 1371 174
rect 1414 182 1415 184
rect 1417 182 1419 184
rect 1414 180 1419 182
rect 1423 217 1428 219
rect 1423 215 1425 217
rect 1427 215 1428 217
rect 1423 213 1428 215
rect 1423 209 1427 213
rect 1423 207 1424 209
rect 1426 207 1427 209
rect 1423 191 1427 207
rect 1502 217 1508 218
rect 1502 215 1503 217
rect 1505 215 1508 217
rect 1502 214 1508 215
rect 1423 189 1428 191
rect 1423 187 1425 189
rect 1427 187 1428 189
rect 1423 182 1428 187
rect 1451 201 1459 203
rect 1471 202 1475 211
rect 1451 199 1452 201
rect 1454 199 1459 201
rect 1451 197 1459 199
rect 1469 201 1484 202
rect 1469 199 1471 201
rect 1473 199 1474 201
rect 1476 199 1478 201
rect 1480 199 1484 201
rect 1469 198 1484 199
rect 1454 194 1459 197
rect 1504 201 1508 214
rect 1504 199 1505 201
rect 1507 199 1508 201
rect 1454 193 1492 194
rect 1454 191 1469 193
rect 1471 191 1492 193
rect 1454 190 1492 191
rect 1504 194 1508 199
rect 1502 192 1508 194
rect 1502 190 1503 192
rect 1505 190 1508 192
rect 1502 185 1508 190
rect 1502 183 1503 185
rect 1505 183 1508 185
rect 1423 180 1425 182
rect 1427 180 1428 182
rect 1423 178 1428 180
rect 1502 181 1508 183
rect 1512 217 1518 218
rect 1512 215 1515 217
rect 1517 215 1518 217
rect 1512 214 1518 215
rect 1592 218 1599 219
rect 1592 217 1596 218
rect 1592 215 1593 217
rect 1595 216 1596 217
rect 1598 216 1599 218
rect 1595 215 1599 216
rect 1512 194 1516 214
rect 1545 209 1549 211
rect 1545 207 1546 209
rect 1548 207 1549 209
rect 1512 192 1518 194
rect 1512 190 1515 192
rect 1517 190 1518 192
rect 1512 188 1518 190
rect 1512 186 1515 188
rect 1517 186 1518 188
rect 1512 185 1518 186
rect 1512 183 1515 185
rect 1517 183 1518 185
rect 1512 181 1518 183
rect 1545 202 1549 207
rect 1592 213 1599 215
rect 1536 201 1551 202
rect 1536 199 1540 201
rect 1542 199 1547 201
rect 1549 199 1551 201
rect 1536 198 1551 199
rect 1561 201 1569 203
rect 1561 199 1566 201
rect 1568 199 1569 201
rect 1561 197 1569 199
rect 1561 196 1566 197
rect 1561 194 1563 196
rect 1565 194 1566 196
rect 1528 190 1566 194
rect 1593 191 1597 213
rect 1602 207 1606 208
rect 1602 205 1603 207
rect 1605 205 1606 207
rect 1602 202 1606 205
rect 1602 201 1623 202
rect 1602 199 1617 201
rect 1619 199 1623 201
rect 1602 198 1623 199
rect 1633 210 1638 212
rect 1633 208 1634 210
rect 1636 208 1638 210
rect 1633 206 1638 208
rect 1592 189 1597 191
rect 1592 187 1593 189
rect 1595 187 1597 189
rect 1592 182 1597 187
rect 1592 180 1593 182
rect 1595 180 1597 182
rect 1602 192 1607 194
rect 1609 192 1623 194
rect 1602 190 1623 192
rect 1602 188 1606 190
rect 1602 186 1603 188
rect 1605 186 1606 188
rect 1602 181 1606 186
rect 1592 178 1597 180
rect 1634 187 1638 206
rect 1657 202 1662 211
rect 1674 215 1686 219
rect 1674 213 1682 215
rect 1684 213 1686 215
rect 1657 201 1671 202
rect 1657 199 1665 201
rect 1667 199 1671 201
rect 1657 198 1671 199
rect 1636 185 1638 187
rect 1634 180 1638 185
rect 1650 193 1663 194
rect 1650 191 1655 193
rect 1657 191 1663 193
rect 1650 190 1663 191
rect 1650 185 1654 190
rect 1682 201 1686 213
rect 1682 199 1683 201
rect 1685 199 1686 201
rect 1682 193 1686 199
rect 1650 183 1651 185
rect 1653 183 1654 185
rect 1650 181 1654 183
rect 1681 191 1686 193
rect 1681 189 1682 191
rect 1684 189 1686 191
rect 1681 184 1686 189
rect 1636 178 1638 180
rect 1625 177 1638 178
rect 1625 175 1627 177
rect 1629 175 1638 177
rect 1625 174 1638 175
rect 1634 173 1638 174
rect 1681 182 1682 184
rect 1684 182 1686 184
rect 1681 180 1686 182
rect 1690 217 1695 219
rect 1690 215 1692 217
rect 1694 215 1695 217
rect 1690 213 1695 215
rect 1690 209 1694 213
rect 1690 207 1691 209
rect 1693 207 1694 209
rect 1690 191 1694 207
rect 1769 217 1775 218
rect 1769 215 1770 217
rect 1772 215 1775 217
rect 1769 214 1775 215
rect 1690 189 1695 191
rect 1690 187 1692 189
rect 1694 187 1695 189
rect 1690 182 1695 187
rect 1718 201 1726 203
rect 1738 202 1742 211
rect 1718 199 1719 201
rect 1721 199 1726 201
rect 1718 197 1726 199
rect 1736 201 1751 202
rect 1736 199 1738 201
rect 1740 199 1741 201
rect 1743 199 1745 201
rect 1747 199 1751 201
rect 1736 198 1751 199
rect 1721 194 1726 197
rect 1771 201 1775 214
rect 1771 199 1772 201
rect 1774 199 1775 201
rect 1721 193 1759 194
rect 1721 191 1736 193
rect 1738 191 1759 193
rect 1721 190 1759 191
rect 1771 194 1775 199
rect 1769 192 1775 194
rect 1769 190 1770 192
rect 1772 190 1775 192
rect 1769 185 1775 190
rect 1769 183 1770 185
rect 1772 183 1775 185
rect 1690 180 1692 182
rect 1694 180 1695 182
rect 1690 178 1695 180
rect 1769 181 1775 183
rect 1779 217 1785 218
rect 1779 215 1782 217
rect 1784 215 1785 217
rect 1779 214 1785 215
rect 1859 218 1866 219
rect 1859 217 1863 218
rect 1859 215 1860 217
rect 1862 216 1863 217
rect 1865 216 1866 218
rect 1862 215 1866 216
rect 1948 217 1972 218
rect 1779 194 1783 214
rect 1812 209 1816 211
rect 1812 207 1813 209
rect 1815 207 1816 209
rect 1779 192 1785 194
rect 1779 190 1782 192
rect 1784 190 1785 192
rect 1779 188 1785 190
rect 1779 186 1782 188
rect 1784 186 1785 188
rect 1779 185 1785 186
rect 1779 183 1782 185
rect 1784 183 1785 185
rect 1779 181 1785 183
rect 1812 202 1816 207
rect 1859 213 1866 215
rect 1948 215 1950 217
rect 1952 215 1972 217
rect 1948 214 1972 215
rect 1803 201 1818 202
rect 1803 199 1807 201
rect 1809 199 1814 201
rect 1816 199 1818 201
rect 1803 198 1818 199
rect 1828 201 1836 203
rect 1828 199 1833 201
rect 1835 199 1836 201
rect 1828 197 1836 199
rect 1828 196 1833 197
rect 1828 194 1830 196
rect 1832 194 1833 196
rect 1795 190 1833 194
rect 1860 191 1864 213
rect 1869 207 1873 208
rect 1869 205 1870 207
rect 1872 205 1873 207
rect 1869 202 1873 205
rect 1869 201 1890 202
rect 1869 199 1884 201
rect 1886 199 1890 201
rect 1869 198 1890 199
rect 1900 210 1905 212
rect 1900 208 1901 210
rect 1903 208 1905 210
rect 1900 206 1905 208
rect 1859 189 1864 191
rect 1859 187 1860 189
rect 1862 187 1864 189
rect 1859 182 1864 187
rect 1859 180 1860 182
rect 1862 180 1864 182
rect 1869 192 1874 194
rect 1876 192 1890 194
rect 1869 190 1890 192
rect 1869 188 1873 190
rect 1869 186 1870 188
rect 1872 186 1873 188
rect 1869 181 1873 186
rect 1859 178 1864 180
rect 1901 187 1905 206
rect 1920 210 1933 211
rect 1920 208 1925 210
rect 1927 208 1933 210
rect 1920 206 1933 208
rect 1920 205 1930 206
rect 1928 204 1930 205
rect 1932 204 1933 206
rect 1903 185 1905 187
rect 1901 180 1905 185
rect 1903 178 1905 180
rect 1892 177 1905 178
rect 1892 175 1894 177
rect 1896 175 1905 177
rect 1892 174 1905 175
rect 1901 173 1905 174
rect 1912 193 1917 195
rect 1912 191 1914 193
rect 1916 191 1917 193
rect 1912 179 1917 191
rect 1928 197 1933 204
rect 1912 173 1924 179
rect 1968 193 1972 214
rect 1968 191 1969 193
rect 1971 191 1972 193
rect 1968 186 1972 191
rect 1956 184 1972 186
rect 1956 182 1958 184
rect 1960 182 1972 184
rect 1956 181 1972 182
rect 1976 217 1981 219
rect 1976 215 1978 217
rect 1980 215 1981 217
rect 1976 213 1981 215
rect 1976 209 1980 213
rect 1976 207 1977 209
rect 1979 207 1980 209
rect 1976 191 1980 207
rect 2055 217 2061 218
rect 2055 215 2056 217
rect 2058 215 2061 217
rect 2055 214 2061 215
rect 1976 189 1981 191
rect 1976 187 1978 189
rect 1980 187 1981 189
rect 1976 182 1981 187
rect 2004 201 2012 203
rect 2024 202 2028 211
rect 2004 199 2005 201
rect 2007 199 2012 201
rect 2004 197 2012 199
rect 2022 201 2037 202
rect 2022 199 2024 201
rect 2026 199 2031 201
rect 2033 199 2037 201
rect 2022 198 2037 199
rect 2007 194 2012 197
rect 2057 201 2061 214
rect 2057 199 2058 201
rect 2060 199 2061 201
rect 2007 193 2045 194
rect 2007 191 2018 193
rect 2020 191 2045 193
rect 2007 190 2045 191
rect 2057 194 2061 199
rect 2055 192 2061 194
rect 2055 190 2056 192
rect 2058 190 2061 192
rect 2055 185 2061 190
rect 2055 183 2056 185
rect 2058 183 2061 185
rect 1976 180 1978 182
rect 1980 180 1981 182
rect 1976 178 1981 180
rect 2055 181 2061 183
rect 2065 217 2071 218
rect 2065 215 2068 217
rect 2070 215 2071 217
rect 2065 214 2071 215
rect 2145 218 2152 219
rect 2145 217 2149 218
rect 2145 215 2146 217
rect 2148 216 2149 217
rect 2151 216 2152 218
rect 2148 215 2152 216
rect 2065 194 2069 214
rect 2098 209 2102 211
rect 2098 207 2099 209
rect 2101 207 2102 209
rect 2065 192 2071 194
rect 2065 190 2068 192
rect 2070 190 2071 192
rect 2065 188 2071 190
rect 2065 186 2068 188
rect 2070 186 2071 188
rect 2065 185 2071 186
rect 2065 183 2068 185
rect 2070 183 2071 185
rect 2065 181 2071 183
rect 2098 202 2102 207
rect 2145 213 2150 215
rect 2089 201 2104 202
rect 2089 199 2093 201
rect 2095 199 2100 201
rect 2102 199 2104 201
rect 2089 198 2104 199
rect 2114 201 2122 203
rect 2114 199 2119 201
rect 2121 199 2122 201
rect 2114 197 2122 199
rect 2114 196 2119 197
rect 2114 194 2116 196
rect 2118 194 2119 196
rect 2081 190 2119 194
rect 2146 191 2150 213
rect 2155 207 2159 211
rect 2155 205 2156 207
rect 2158 205 2159 207
rect 2155 202 2159 205
rect 2155 201 2176 202
rect 2155 199 2170 201
rect 2172 199 2176 201
rect 2155 198 2176 199
rect 2186 210 2191 212
rect 2186 208 2187 210
rect 2189 208 2191 210
rect 2186 206 2191 208
rect 2145 189 2150 191
rect 2145 187 2146 189
rect 2148 187 2150 189
rect 2145 182 2150 187
rect 2145 180 2146 182
rect 2148 180 2150 182
rect 2155 192 2160 194
rect 2162 192 2176 194
rect 2155 190 2176 192
rect 2155 188 2159 190
rect 2155 186 2156 188
rect 2158 186 2159 188
rect 2155 181 2159 186
rect 2145 178 2150 180
rect 2187 187 2191 206
rect 2255 217 2259 219
rect 2254 215 2259 217
rect 2254 213 2255 215
rect 2257 213 2259 215
rect 2254 211 2259 213
rect 2206 209 2219 210
rect 2206 207 2210 209
rect 2212 207 2219 209
rect 2206 206 2219 207
rect 2213 201 2219 206
rect 2213 199 2214 201
rect 2216 199 2219 201
rect 2213 197 2219 199
rect 2239 196 2243 203
rect 2239 195 2241 196
rect 2231 194 2241 195
rect 2231 193 2243 194
rect 2231 191 2236 193
rect 2238 191 2243 193
rect 2231 189 2243 191
rect 2189 185 2191 187
rect 2187 180 2191 185
rect 2189 178 2191 180
rect 2178 177 2191 178
rect 2178 175 2180 177
rect 2182 175 2191 177
rect 2178 174 2191 175
rect 2187 173 2191 174
rect 2199 182 2212 186
rect 2199 181 2204 182
rect 2199 179 2201 181
rect 2203 179 2204 181
rect 2199 173 2204 179
rect 2255 178 2259 211
rect 2323 217 2327 219
rect 2322 215 2327 217
rect 2322 213 2323 215
rect 2325 213 2327 215
rect 2322 211 2327 213
rect 2274 209 2287 210
rect 2274 207 2276 209
rect 2278 207 2287 209
rect 2274 206 2287 207
rect 2281 201 2287 206
rect 2281 199 2282 201
rect 2284 199 2287 201
rect 2281 197 2287 199
rect 2307 196 2311 203
rect 2307 195 2309 196
rect 2299 194 2309 195
rect 2299 192 2300 194
rect 2302 192 2311 194
rect 2299 189 2311 192
rect 2246 177 2259 178
rect 2246 175 2255 177
rect 2257 175 2259 177
rect 2246 174 2259 175
rect 2267 182 2280 186
rect 2267 181 2272 182
rect 2267 179 2269 181
rect 2271 179 2272 181
rect 2267 173 2272 179
rect 2323 178 2327 211
rect 2314 177 2327 178
rect 2314 175 2323 177
rect 2325 175 2327 177
rect 2314 174 2327 175
rect 4 167 306 168
rect 4 165 39 167
rect 41 165 79 167
rect 81 165 298 167
rect 300 165 306 167
rect 4 155 306 165
rect 4 153 39 155
rect 41 153 79 155
rect 81 153 298 155
rect 300 153 306 155
rect 4 152 306 153
rect 311 167 573 168
rect 311 165 346 167
rect 348 165 565 167
rect 567 165 573 167
rect 311 155 573 165
rect 311 153 346 155
rect 348 153 565 155
rect 567 153 573 155
rect 311 152 573 153
rect 578 167 840 168
rect 578 165 613 167
rect 615 165 832 167
rect 834 165 840 167
rect 578 155 840 165
rect 578 153 613 155
rect 615 153 832 155
rect 834 153 840 155
rect 578 152 840 153
rect 845 167 1107 168
rect 845 165 880 167
rect 882 165 1099 167
rect 1101 165 1107 167
rect 845 155 1107 165
rect 845 153 880 155
rect 882 153 1099 155
rect 1101 153 1107 155
rect 845 152 1107 153
rect 1112 167 1374 168
rect 1112 165 1147 167
rect 1149 165 1366 167
rect 1368 165 1374 167
rect 1112 155 1374 165
rect 1112 153 1147 155
rect 1149 153 1366 155
rect 1368 153 1374 155
rect 1112 152 1374 153
rect 1379 167 1641 168
rect 1379 165 1414 167
rect 1416 165 1633 167
rect 1635 165 1641 167
rect 1379 155 1641 165
rect 1379 153 1414 155
rect 1416 153 1633 155
rect 1635 153 1641 155
rect 1379 152 1641 153
rect 1646 167 2331 168
rect 1646 165 1681 167
rect 1683 165 1900 167
rect 1902 165 1948 167
rect 1950 165 2186 167
rect 2188 165 2320 167
rect 2322 165 2331 167
rect 1646 155 2331 165
rect 1646 153 1681 155
rect 1683 153 1900 155
rect 1902 153 1948 155
rect 1950 153 2186 155
rect 2188 153 2331 155
rect 1646 152 2331 153
rect 8 132 12 139
rect 39 141 44 143
rect 39 139 40 141
rect 42 139 44 141
rect 8 130 9 132
rect 11 130 12 132
rect 8 129 21 130
rect 8 127 13 129
rect 15 127 21 129
rect 8 126 21 127
rect 15 121 29 122
rect 15 119 23 121
rect 25 119 29 121
rect 15 118 29 119
rect 39 133 44 139
rect 39 131 40 133
rect 42 131 44 133
rect 39 129 44 131
rect 39 127 41 129
rect 43 127 44 129
rect 39 125 44 127
rect 48 130 52 139
rect 299 146 303 147
rect 290 142 303 146
rect 88 140 93 142
rect 79 138 84 140
rect 48 129 61 130
rect 48 127 53 129
rect 55 127 61 129
rect 48 126 61 127
rect 15 109 20 118
rect 40 107 44 125
rect 55 121 69 122
rect 55 119 63 121
rect 65 119 69 121
rect 55 118 69 119
rect 79 136 80 138
rect 82 136 84 138
rect 79 131 84 136
rect 79 129 80 131
rect 82 129 84 131
rect 79 127 84 129
rect 55 116 60 118
rect 55 114 57 116
rect 59 114 60 116
rect 55 109 60 114
rect 80 121 84 127
rect 80 119 81 121
rect 83 119 84 121
rect 32 105 40 107
rect 42 105 44 107
rect 80 107 84 119
rect 32 101 44 105
rect 72 105 80 107
rect 82 105 84 107
rect 72 101 84 105
rect 88 138 90 140
rect 92 138 93 140
rect 88 133 93 138
rect 88 131 90 133
rect 92 131 93 133
rect 88 129 93 131
rect 88 113 92 129
rect 119 129 157 130
rect 119 127 138 129
rect 140 127 157 129
rect 119 126 157 127
rect 119 123 124 126
rect 116 121 124 123
rect 116 119 117 121
rect 119 119 124 121
rect 116 117 124 119
rect 134 121 149 122
rect 134 119 136 121
rect 138 119 140 121
rect 142 119 143 121
rect 145 119 149 121
rect 134 118 149 119
rect 88 111 89 113
rect 91 111 92 113
rect 88 107 92 111
rect 88 105 93 107
rect 136 109 140 118
rect 167 137 173 139
rect 167 135 168 137
rect 170 135 173 137
rect 167 130 173 135
rect 167 128 168 130
rect 170 128 173 130
rect 167 126 173 128
rect 169 121 173 126
rect 169 119 170 121
rect 172 119 173 121
rect 169 106 173 119
rect 88 103 90 105
rect 92 103 93 105
rect 88 101 93 103
rect 167 105 173 106
rect 167 103 168 105
rect 170 103 173 105
rect 167 102 173 103
rect 177 137 183 139
rect 257 140 262 142
rect 257 138 258 140
rect 260 138 262 140
rect 177 135 180 137
rect 182 135 183 137
rect 177 134 183 135
rect 177 132 180 134
rect 182 132 183 134
rect 177 130 183 132
rect 177 128 180 130
rect 182 128 183 130
rect 177 126 183 128
rect 177 106 181 126
rect 193 129 231 130
rect 193 127 228 129
rect 230 127 231 129
rect 193 126 231 127
rect 226 123 231 126
rect 201 121 216 122
rect 201 119 205 121
rect 207 119 212 121
rect 214 119 216 121
rect 201 118 216 119
rect 226 121 234 123
rect 226 119 231 121
rect 233 119 234 121
rect 210 113 214 118
rect 226 117 234 119
rect 257 133 262 138
rect 257 131 258 133
rect 260 131 262 133
rect 257 129 262 131
rect 210 111 211 113
rect 213 111 214 113
rect 210 109 214 111
rect 177 105 183 106
rect 177 103 180 105
rect 182 103 183 105
rect 177 102 183 103
rect 258 107 262 129
rect 267 138 271 139
rect 267 136 268 138
rect 270 136 271 138
rect 267 130 271 136
rect 267 128 288 130
rect 267 126 272 128
rect 274 126 288 128
rect 267 121 288 122
rect 267 119 268 121
rect 270 119 282 121
rect 284 119 288 121
rect 267 118 288 119
rect 301 140 303 142
rect 299 135 303 140
rect 301 133 303 135
rect 267 114 271 118
rect 299 117 303 133
rect 315 130 319 139
rect 566 146 570 147
rect 557 142 570 146
rect 355 140 360 142
rect 346 138 351 140
rect 315 129 328 130
rect 315 127 320 129
rect 322 127 328 129
rect 315 126 328 127
rect 299 115 300 117
rect 302 115 303 117
rect 299 114 303 115
rect 298 112 303 114
rect 298 110 299 112
rect 301 110 303 112
rect 298 108 303 110
rect 322 121 336 122
rect 322 119 330 121
rect 332 119 336 121
rect 322 118 336 119
rect 346 136 347 138
rect 349 136 351 138
rect 346 131 351 136
rect 346 129 347 131
rect 349 129 351 131
rect 346 127 351 129
rect 322 116 327 118
rect 322 114 324 116
rect 326 114 327 116
rect 322 109 327 114
rect 347 121 351 127
rect 347 119 348 121
rect 350 119 351 121
rect 257 105 264 107
rect 347 107 351 119
rect 257 103 258 105
rect 260 104 264 105
rect 260 103 261 104
rect 257 102 261 103
rect 263 102 264 104
rect 339 105 347 107
rect 349 105 351 107
rect 257 101 264 102
rect 339 101 351 105
rect 355 138 357 140
rect 359 138 360 140
rect 355 133 360 138
rect 355 131 357 133
rect 359 131 360 133
rect 355 129 360 131
rect 355 113 359 129
rect 386 129 424 130
rect 386 127 405 129
rect 407 127 424 129
rect 386 126 424 127
rect 386 123 391 126
rect 383 121 391 123
rect 383 119 384 121
rect 386 119 391 121
rect 383 117 391 119
rect 401 121 416 122
rect 401 119 403 121
rect 405 119 407 121
rect 409 119 410 121
rect 412 119 416 121
rect 401 118 416 119
rect 355 111 356 113
rect 358 111 359 113
rect 355 107 359 111
rect 355 105 360 107
rect 403 109 407 118
rect 434 137 440 139
rect 434 135 435 137
rect 437 135 440 137
rect 434 130 440 135
rect 434 128 435 130
rect 437 128 440 130
rect 434 126 440 128
rect 436 121 440 126
rect 436 119 437 121
rect 439 119 440 121
rect 436 106 440 119
rect 355 103 357 105
rect 359 103 360 105
rect 355 101 360 103
rect 434 105 440 106
rect 434 103 435 105
rect 437 103 440 105
rect 434 102 440 103
rect 444 137 450 139
rect 524 140 529 142
rect 524 138 525 140
rect 527 138 529 140
rect 444 135 447 137
rect 449 135 450 137
rect 444 134 450 135
rect 444 132 447 134
rect 449 132 450 134
rect 444 130 450 132
rect 444 128 447 130
rect 449 128 450 130
rect 444 126 450 128
rect 444 106 448 126
rect 460 129 498 130
rect 460 127 495 129
rect 497 127 498 129
rect 460 126 498 127
rect 493 123 498 126
rect 468 121 483 122
rect 468 119 472 121
rect 474 119 479 121
rect 481 119 483 121
rect 468 118 483 119
rect 493 121 501 123
rect 493 119 498 121
rect 500 119 501 121
rect 477 113 481 118
rect 493 117 501 119
rect 524 133 529 138
rect 524 131 525 133
rect 527 131 529 133
rect 524 129 529 131
rect 477 111 478 113
rect 480 111 481 113
rect 477 109 481 111
rect 444 105 450 106
rect 444 103 447 105
rect 449 103 450 105
rect 444 102 450 103
rect 525 107 529 129
rect 534 138 538 139
rect 534 136 535 138
rect 537 136 538 138
rect 534 130 538 136
rect 534 128 555 130
rect 534 126 539 128
rect 541 126 555 128
rect 534 121 555 122
rect 534 119 535 121
rect 537 119 549 121
rect 551 119 555 121
rect 534 118 555 119
rect 568 140 570 142
rect 566 135 570 140
rect 568 133 570 135
rect 534 114 538 118
rect 566 117 570 133
rect 582 130 586 139
rect 833 146 837 147
rect 824 142 837 146
rect 622 140 627 142
rect 613 138 618 140
rect 582 129 595 130
rect 582 127 587 129
rect 589 127 595 129
rect 582 126 595 127
rect 566 115 567 117
rect 569 115 570 117
rect 566 114 570 115
rect 565 112 570 114
rect 565 110 566 112
rect 568 110 570 112
rect 565 108 570 110
rect 589 121 603 122
rect 589 119 597 121
rect 599 119 603 121
rect 589 118 603 119
rect 613 136 614 138
rect 616 136 618 138
rect 613 131 618 136
rect 613 129 614 131
rect 616 129 618 131
rect 613 127 618 129
rect 589 116 594 118
rect 589 114 591 116
rect 593 114 594 116
rect 589 109 594 114
rect 614 121 618 127
rect 614 119 615 121
rect 617 119 618 121
rect 524 105 531 107
rect 614 107 618 119
rect 524 103 525 105
rect 527 104 531 105
rect 527 103 528 104
rect 524 102 528 103
rect 530 102 531 104
rect 606 105 614 107
rect 616 105 618 107
rect 524 101 531 102
rect 606 101 618 105
rect 622 138 624 140
rect 626 138 627 140
rect 622 133 627 138
rect 622 131 624 133
rect 626 131 627 133
rect 622 129 627 131
rect 622 113 626 129
rect 653 129 691 130
rect 653 127 672 129
rect 674 127 691 129
rect 653 126 691 127
rect 653 123 658 126
rect 650 121 658 123
rect 650 119 651 121
rect 653 119 658 121
rect 650 117 658 119
rect 668 121 683 122
rect 668 119 670 121
rect 672 119 674 121
rect 676 119 677 121
rect 679 119 683 121
rect 668 118 683 119
rect 622 111 623 113
rect 625 111 626 113
rect 622 107 626 111
rect 622 105 627 107
rect 670 109 674 118
rect 701 137 707 139
rect 701 135 702 137
rect 704 135 707 137
rect 701 130 707 135
rect 701 128 702 130
rect 704 128 707 130
rect 701 126 707 128
rect 703 121 707 126
rect 703 119 704 121
rect 706 119 707 121
rect 703 106 707 119
rect 622 103 624 105
rect 626 103 627 105
rect 622 101 627 103
rect 701 105 707 106
rect 701 103 702 105
rect 704 103 707 105
rect 701 102 707 103
rect 711 137 717 139
rect 791 140 796 142
rect 791 138 792 140
rect 794 138 796 140
rect 711 135 714 137
rect 716 135 717 137
rect 711 134 717 135
rect 711 132 714 134
rect 716 132 717 134
rect 711 130 717 132
rect 711 128 714 130
rect 716 128 717 130
rect 711 126 717 128
rect 711 106 715 126
rect 727 129 765 130
rect 727 127 762 129
rect 764 127 765 129
rect 727 126 765 127
rect 760 123 765 126
rect 735 121 750 122
rect 735 119 739 121
rect 741 119 746 121
rect 748 119 750 121
rect 735 118 750 119
rect 760 121 768 123
rect 760 119 765 121
rect 767 119 768 121
rect 744 113 748 118
rect 760 117 768 119
rect 791 133 796 138
rect 791 131 792 133
rect 794 131 796 133
rect 791 129 796 131
rect 744 111 745 113
rect 747 111 748 113
rect 744 109 748 111
rect 711 105 717 106
rect 711 103 714 105
rect 716 103 717 105
rect 711 102 717 103
rect 792 107 796 129
rect 801 138 805 139
rect 801 136 802 138
rect 804 136 805 138
rect 801 130 805 136
rect 801 128 822 130
rect 801 126 806 128
rect 808 126 822 128
rect 801 121 822 122
rect 801 119 802 121
rect 804 119 816 121
rect 818 119 822 121
rect 801 118 822 119
rect 835 140 837 142
rect 833 135 837 140
rect 835 133 837 135
rect 801 114 805 118
rect 833 117 837 133
rect 849 130 853 139
rect 1100 146 1104 147
rect 1091 142 1104 146
rect 889 140 894 142
rect 880 138 885 140
rect 849 129 862 130
rect 849 127 854 129
rect 856 127 862 129
rect 849 126 862 127
rect 833 115 834 117
rect 836 115 837 117
rect 833 114 837 115
rect 832 112 837 114
rect 832 110 833 112
rect 835 110 837 112
rect 832 108 837 110
rect 856 121 870 122
rect 856 119 864 121
rect 866 119 870 121
rect 856 118 870 119
rect 880 136 881 138
rect 883 136 885 138
rect 880 131 885 136
rect 880 129 881 131
rect 883 129 885 131
rect 880 127 885 129
rect 856 116 861 118
rect 856 114 858 116
rect 860 114 861 116
rect 856 109 861 114
rect 881 121 885 127
rect 881 119 882 121
rect 884 119 885 121
rect 791 105 798 107
rect 881 107 885 119
rect 791 103 792 105
rect 794 104 798 105
rect 794 103 795 104
rect 791 102 795 103
rect 797 102 798 104
rect 873 105 881 107
rect 883 105 885 107
rect 791 101 798 102
rect 873 101 885 105
rect 889 138 891 140
rect 893 138 894 140
rect 889 133 894 138
rect 889 131 891 133
rect 893 131 894 133
rect 889 129 894 131
rect 889 113 893 129
rect 920 129 958 130
rect 920 127 939 129
rect 941 127 958 129
rect 920 126 958 127
rect 920 123 925 126
rect 917 121 925 123
rect 917 119 918 121
rect 920 119 925 121
rect 917 117 925 119
rect 935 121 950 122
rect 935 119 937 121
rect 939 119 941 121
rect 943 119 944 121
rect 946 119 950 121
rect 935 118 950 119
rect 889 111 890 113
rect 892 111 893 113
rect 889 107 893 111
rect 889 105 894 107
rect 937 109 941 118
rect 968 137 974 139
rect 968 135 969 137
rect 971 135 974 137
rect 968 130 974 135
rect 968 128 969 130
rect 971 128 974 130
rect 968 126 974 128
rect 970 121 974 126
rect 970 119 971 121
rect 973 119 974 121
rect 970 106 974 119
rect 889 103 891 105
rect 893 103 894 105
rect 889 101 894 103
rect 968 105 974 106
rect 968 103 969 105
rect 971 103 974 105
rect 968 102 974 103
rect 978 137 984 139
rect 1058 140 1063 142
rect 1058 138 1059 140
rect 1061 138 1063 140
rect 978 135 981 137
rect 983 135 984 137
rect 978 134 984 135
rect 978 132 981 134
rect 983 132 984 134
rect 978 130 984 132
rect 978 128 981 130
rect 983 128 984 130
rect 978 126 984 128
rect 978 106 982 126
rect 994 129 1032 130
rect 994 127 1029 129
rect 1031 127 1032 129
rect 994 126 1032 127
rect 1027 123 1032 126
rect 1002 121 1017 122
rect 1002 119 1006 121
rect 1008 119 1013 121
rect 1015 119 1017 121
rect 1002 118 1017 119
rect 1027 121 1035 123
rect 1027 119 1032 121
rect 1034 119 1035 121
rect 1011 113 1015 118
rect 1027 117 1035 119
rect 1058 133 1063 138
rect 1058 131 1059 133
rect 1061 131 1063 133
rect 1058 129 1063 131
rect 1011 111 1012 113
rect 1014 111 1015 113
rect 1011 109 1015 111
rect 978 105 984 106
rect 978 103 981 105
rect 983 103 984 105
rect 978 102 984 103
rect 1059 107 1063 129
rect 1068 138 1072 139
rect 1068 136 1069 138
rect 1071 136 1072 138
rect 1068 130 1072 136
rect 1068 128 1089 130
rect 1068 126 1073 128
rect 1075 126 1089 128
rect 1068 121 1089 122
rect 1068 119 1069 121
rect 1071 119 1083 121
rect 1085 119 1089 121
rect 1068 118 1089 119
rect 1102 140 1104 142
rect 1100 135 1104 140
rect 1102 133 1104 135
rect 1068 114 1072 118
rect 1100 117 1104 133
rect 1116 130 1120 139
rect 1367 146 1371 147
rect 1358 142 1371 146
rect 1156 140 1161 142
rect 1147 138 1152 140
rect 1116 129 1129 130
rect 1116 127 1121 129
rect 1123 127 1129 129
rect 1116 126 1129 127
rect 1100 115 1101 117
rect 1103 115 1104 117
rect 1100 114 1104 115
rect 1099 112 1104 114
rect 1099 110 1100 112
rect 1102 110 1104 112
rect 1099 108 1104 110
rect 1123 121 1137 122
rect 1123 119 1131 121
rect 1133 119 1137 121
rect 1123 118 1137 119
rect 1147 136 1148 138
rect 1150 136 1152 138
rect 1147 131 1152 136
rect 1147 129 1148 131
rect 1150 129 1152 131
rect 1147 127 1152 129
rect 1123 116 1128 118
rect 1123 114 1125 116
rect 1127 114 1128 116
rect 1123 109 1128 114
rect 1148 121 1152 127
rect 1148 119 1149 121
rect 1151 119 1152 121
rect 1058 105 1065 107
rect 1148 107 1152 119
rect 1058 103 1059 105
rect 1061 104 1065 105
rect 1061 103 1062 104
rect 1058 102 1062 103
rect 1064 102 1065 104
rect 1140 105 1148 107
rect 1150 105 1152 107
rect 1058 101 1065 102
rect 1140 101 1152 105
rect 1156 138 1158 140
rect 1160 138 1161 140
rect 1156 133 1161 138
rect 1156 131 1158 133
rect 1160 131 1161 133
rect 1156 129 1161 131
rect 1156 113 1160 129
rect 1187 129 1225 130
rect 1187 127 1206 129
rect 1208 127 1225 129
rect 1187 126 1225 127
rect 1187 123 1192 126
rect 1184 121 1192 123
rect 1184 119 1185 121
rect 1187 119 1192 121
rect 1184 117 1192 119
rect 1202 121 1217 122
rect 1202 119 1204 121
rect 1206 119 1208 121
rect 1210 119 1211 121
rect 1213 119 1217 121
rect 1202 118 1217 119
rect 1156 111 1157 113
rect 1159 111 1160 113
rect 1156 107 1160 111
rect 1156 105 1161 107
rect 1204 109 1208 118
rect 1235 137 1241 139
rect 1235 135 1236 137
rect 1238 135 1241 137
rect 1235 130 1241 135
rect 1235 128 1236 130
rect 1238 128 1241 130
rect 1235 126 1241 128
rect 1237 121 1241 126
rect 1237 119 1238 121
rect 1240 119 1241 121
rect 1237 106 1241 119
rect 1156 103 1158 105
rect 1160 103 1161 105
rect 1156 101 1161 103
rect 1235 105 1241 106
rect 1235 103 1236 105
rect 1238 103 1241 105
rect 1235 102 1241 103
rect 1245 137 1251 139
rect 1325 140 1330 142
rect 1325 138 1326 140
rect 1328 138 1330 140
rect 1245 135 1248 137
rect 1250 135 1251 137
rect 1245 134 1251 135
rect 1245 132 1248 134
rect 1250 132 1251 134
rect 1245 130 1251 132
rect 1245 128 1248 130
rect 1250 128 1251 130
rect 1245 126 1251 128
rect 1245 106 1249 126
rect 1261 129 1299 130
rect 1261 127 1296 129
rect 1298 127 1299 129
rect 1261 126 1299 127
rect 1294 123 1299 126
rect 1269 121 1284 122
rect 1269 119 1273 121
rect 1275 119 1280 121
rect 1282 119 1284 121
rect 1269 118 1284 119
rect 1294 121 1302 123
rect 1294 119 1299 121
rect 1301 119 1302 121
rect 1278 113 1282 118
rect 1294 117 1302 119
rect 1325 133 1330 138
rect 1325 131 1326 133
rect 1328 131 1330 133
rect 1325 129 1330 131
rect 1278 111 1279 113
rect 1281 111 1282 113
rect 1278 109 1282 111
rect 1245 105 1251 106
rect 1245 103 1248 105
rect 1250 103 1251 105
rect 1245 102 1251 103
rect 1326 107 1330 129
rect 1335 138 1339 139
rect 1335 136 1336 138
rect 1338 136 1339 138
rect 1335 130 1339 136
rect 1335 128 1356 130
rect 1335 126 1340 128
rect 1342 126 1356 128
rect 1335 121 1356 122
rect 1335 119 1336 121
rect 1338 119 1350 121
rect 1352 119 1356 121
rect 1335 118 1356 119
rect 1369 140 1371 142
rect 1367 135 1371 140
rect 1369 133 1371 135
rect 1335 114 1339 118
rect 1367 117 1371 133
rect 1383 130 1387 139
rect 1634 146 1638 147
rect 1625 142 1638 146
rect 1423 140 1428 142
rect 1414 138 1419 140
rect 1383 129 1396 130
rect 1383 127 1388 129
rect 1390 127 1396 129
rect 1383 126 1396 127
rect 1367 115 1368 117
rect 1370 115 1371 117
rect 1367 114 1371 115
rect 1366 112 1371 114
rect 1366 110 1367 112
rect 1369 110 1371 112
rect 1366 108 1371 110
rect 1390 121 1404 122
rect 1390 119 1398 121
rect 1400 119 1404 121
rect 1390 118 1404 119
rect 1414 136 1415 138
rect 1417 136 1419 138
rect 1414 131 1419 136
rect 1414 129 1415 131
rect 1417 129 1419 131
rect 1414 127 1419 129
rect 1390 116 1395 118
rect 1390 114 1392 116
rect 1394 114 1395 116
rect 1390 109 1395 114
rect 1415 121 1419 127
rect 1415 119 1416 121
rect 1418 119 1419 121
rect 1325 105 1332 107
rect 1415 107 1419 119
rect 1325 103 1326 105
rect 1328 104 1332 105
rect 1328 103 1329 104
rect 1325 102 1329 103
rect 1331 102 1332 104
rect 1407 105 1415 107
rect 1417 105 1419 107
rect 1325 101 1332 102
rect 1407 101 1419 105
rect 1423 138 1425 140
rect 1427 138 1428 140
rect 1423 133 1428 138
rect 1423 131 1425 133
rect 1427 131 1428 133
rect 1423 129 1428 131
rect 1423 113 1427 129
rect 1454 129 1492 130
rect 1454 127 1473 129
rect 1475 127 1492 129
rect 1454 126 1492 127
rect 1454 123 1459 126
rect 1451 121 1459 123
rect 1451 119 1452 121
rect 1454 119 1459 121
rect 1451 117 1459 119
rect 1469 121 1484 122
rect 1469 119 1471 121
rect 1473 119 1475 121
rect 1477 119 1478 121
rect 1480 119 1484 121
rect 1469 118 1484 119
rect 1423 111 1424 113
rect 1426 111 1427 113
rect 1423 107 1427 111
rect 1423 105 1428 107
rect 1471 109 1475 118
rect 1502 137 1508 139
rect 1502 135 1503 137
rect 1505 135 1508 137
rect 1502 130 1508 135
rect 1502 128 1503 130
rect 1505 128 1508 130
rect 1502 126 1508 128
rect 1504 121 1508 126
rect 1504 119 1505 121
rect 1507 119 1508 121
rect 1504 106 1508 119
rect 1423 103 1425 105
rect 1427 103 1428 105
rect 1423 101 1428 103
rect 1502 105 1508 106
rect 1502 103 1503 105
rect 1505 103 1508 105
rect 1502 102 1508 103
rect 1512 137 1518 139
rect 1592 140 1597 142
rect 1592 138 1593 140
rect 1595 138 1597 140
rect 1512 135 1515 137
rect 1517 135 1518 137
rect 1512 134 1518 135
rect 1512 132 1515 134
rect 1517 132 1518 134
rect 1512 130 1518 132
rect 1512 128 1515 130
rect 1517 128 1518 130
rect 1512 126 1518 128
rect 1512 106 1516 126
rect 1528 129 1566 130
rect 1528 127 1563 129
rect 1565 127 1566 129
rect 1528 126 1566 127
rect 1561 123 1566 126
rect 1536 121 1551 122
rect 1536 119 1540 121
rect 1542 119 1547 121
rect 1549 119 1551 121
rect 1536 118 1551 119
rect 1561 121 1569 123
rect 1561 119 1566 121
rect 1568 119 1569 121
rect 1545 113 1549 118
rect 1561 117 1569 119
rect 1592 133 1597 138
rect 1592 131 1593 133
rect 1595 131 1597 133
rect 1592 129 1597 131
rect 1545 111 1546 113
rect 1548 111 1549 113
rect 1545 109 1549 111
rect 1512 105 1518 106
rect 1512 103 1515 105
rect 1517 103 1518 105
rect 1512 102 1518 103
rect 1593 107 1597 129
rect 1602 138 1606 139
rect 1602 136 1603 138
rect 1605 136 1606 138
rect 1602 130 1606 136
rect 1602 128 1623 130
rect 1602 126 1607 128
rect 1609 126 1623 128
rect 1602 121 1623 122
rect 1602 119 1603 121
rect 1605 119 1617 121
rect 1619 119 1623 121
rect 1602 118 1623 119
rect 1636 140 1638 142
rect 1634 135 1638 140
rect 1636 133 1638 135
rect 1602 114 1606 118
rect 1634 117 1638 133
rect 1650 130 1654 139
rect 1901 146 1905 147
rect 1892 142 1905 146
rect 1690 140 1695 142
rect 1681 138 1686 140
rect 1650 129 1663 130
rect 1650 127 1655 129
rect 1657 127 1663 129
rect 1650 126 1663 127
rect 1634 115 1635 117
rect 1637 115 1638 117
rect 1634 114 1638 115
rect 1633 112 1638 114
rect 1633 110 1634 112
rect 1636 110 1638 112
rect 1633 108 1638 110
rect 1657 121 1671 122
rect 1657 119 1665 121
rect 1667 119 1671 121
rect 1657 118 1671 119
rect 1681 136 1682 138
rect 1684 136 1686 138
rect 1681 131 1686 136
rect 1681 129 1682 131
rect 1684 129 1686 131
rect 1681 127 1686 129
rect 1657 116 1662 118
rect 1657 114 1659 116
rect 1661 114 1662 116
rect 1657 109 1662 114
rect 1682 121 1686 127
rect 1682 119 1683 121
rect 1685 119 1686 121
rect 1592 105 1599 107
rect 1682 107 1686 119
rect 1592 103 1593 105
rect 1595 104 1599 105
rect 1595 103 1596 104
rect 1592 102 1596 103
rect 1598 102 1599 104
rect 1674 105 1682 107
rect 1684 105 1686 107
rect 1592 101 1599 102
rect 1674 101 1686 105
rect 1690 138 1692 140
rect 1694 138 1695 140
rect 1690 133 1695 138
rect 1690 131 1692 133
rect 1694 131 1695 133
rect 1690 129 1695 131
rect 1690 113 1694 129
rect 1721 129 1759 130
rect 1721 127 1740 129
rect 1742 127 1759 129
rect 1721 126 1759 127
rect 1721 123 1726 126
rect 1718 121 1726 123
rect 1718 119 1719 121
rect 1721 119 1726 121
rect 1718 117 1726 119
rect 1736 121 1751 122
rect 1736 119 1738 121
rect 1740 119 1742 121
rect 1744 119 1745 121
rect 1747 119 1751 121
rect 1736 118 1751 119
rect 1690 111 1691 113
rect 1693 111 1694 113
rect 1690 107 1694 111
rect 1690 105 1695 107
rect 1738 109 1742 118
rect 1769 137 1775 139
rect 1769 135 1770 137
rect 1772 135 1775 137
rect 1769 130 1775 135
rect 1769 128 1770 130
rect 1772 128 1775 130
rect 1769 126 1775 128
rect 1771 121 1775 126
rect 1771 119 1772 121
rect 1774 119 1775 121
rect 1771 106 1775 119
rect 1690 103 1692 105
rect 1694 103 1695 105
rect 1690 101 1695 103
rect 1769 105 1775 106
rect 1769 103 1770 105
rect 1772 103 1775 105
rect 1769 102 1775 103
rect 1779 137 1785 139
rect 1859 140 1864 142
rect 1859 138 1860 140
rect 1862 138 1864 140
rect 1779 135 1782 137
rect 1784 135 1785 137
rect 1779 134 1785 135
rect 1779 132 1782 134
rect 1784 132 1785 134
rect 1779 130 1785 132
rect 1779 128 1782 130
rect 1784 128 1785 130
rect 1779 126 1785 128
rect 1779 106 1783 126
rect 1795 129 1833 130
rect 1795 127 1830 129
rect 1832 127 1833 129
rect 1795 126 1833 127
rect 1828 123 1833 126
rect 1803 121 1818 122
rect 1803 119 1807 121
rect 1809 119 1814 121
rect 1816 119 1818 121
rect 1803 118 1818 119
rect 1828 121 1836 123
rect 1828 119 1833 121
rect 1835 119 1836 121
rect 1812 113 1816 118
rect 1828 117 1836 119
rect 1859 133 1864 138
rect 1859 131 1860 133
rect 1862 131 1864 133
rect 1859 129 1864 131
rect 1812 111 1813 113
rect 1815 111 1816 113
rect 1812 109 1816 111
rect 1779 105 1785 106
rect 1779 103 1782 105
rect 1784 103 1785 105
rect 1779 102 1785 103
rect 1860 113 1864 129
rect 1869 138 1873 139
rect 1869 136 1870 138
rect 1872 136 1873 138
rect 1869 130 1873 136
rect 1869 128 1890 130
rect 1869 126 1874 128
rect 1876 126 1890 128
rect 1869 121 1890 122
rect 1869 119 1870 121
rect 1872 119 1884 121
rect 1886 119 1890 121
rect 1869 118 1890 119
rect 1903 140 1905 142
rect 1901 135 1905 140
rect 1903 133 1905 135
rect 1869 114 1873 118
rect 1901 117 1905 133
rect 1912 141 1924 147
rect 1912 129 1917 141
rect 2187 146 2191 147
rect 2178 142 2191 146
rect 1976 140 1981 142
rect 1912 127 1914 129
rect 1916 127 1917 129
rect 1912 125 1917 127
rect 1901 115 1902 117
rect 1904 115 1905 117
rect 1901 114 1905 115
rect 1860 111 1861 113
rect 1863 111 1864 113
rect 1860 107 1864 111
rect 1900 112 1905 114
rect 1900 110 1901 112
rect 1903 110 1905 112
rect 1900 108 1905 110
rect 1928 116 1933 123
rect 1956 138 1972 139
rect 1956 136 1958 138
rect 1960 136 1972 138
rect 1956 134 1972 136
rect 1968 129 1972 134
rect 1968 127 1969 129
rect 1971 127 1972 129
rect 1928 115 1930 116
rect 1920 114 1930 115
rect 1932 114 1933 116
rect 1920 112 1933 114
rect 1920 110 1925 112
rect 1927 110 1933 112
rect 1920 109 1933 110
rect 1859 105 1866 107
rect 1968 106 1972 127
rect 1859 103 1860 105
rect 1862 103 1866 105
rect 1859 101 1866 103
rect 1948 105 1972 106
rect 1948 103 1950 105
rect 1952 103 1972 105
rect 1948 102 1972 103
rect 1976 138 1978 140
rect 1980 138 1981 140
rect 1976 133 1981 138
rect 1976 131 1978 133
rect 1980 131 1981 133
rect 1976 129 1981 131
rect 1976 113 1980 129
rect 2007 129 2045 130
rect 2007 127 2018 129
rect 2020 127 2045 129
rect 2007 126 2045 127
rect 2007 123 2012 126
rect 2004 121 2012 123
rect 2004 119 2005 121
rect 2007 119 2012 121
rect 2004 117 2012 119
rect 2022 121 2037 122
rect 2022 119 2024 121
rect 2026 119 2031 121
rect 2033 119 2037 121
rect 2022 118 2037 119
rect 1976 111 1977 113
rect 1979 111 1980 113
rect 1976 107 1980 111
rect 1976 105 1981 107
rect 2024 109 2028 118
rect 2055 137 2061 139
rect 2055 135 2056 137
rect 2058 135 2061 137
rect 2055 130 2061 135
rect 2055 128 2056 130
rect 2058 128 2061 130
rect 2055 126 2061 128
rect 2057 121 2061 126
rect 2057 119 2058 121
rect 2060 119 2061 121
rect 2057 106 2061 119
rect 1976 103 1978 105
rect 1980 103 1981 105
rect 1976 101 1981 103
rect 2055 105 2061 106
rect 2055 103 2056 105
rect 2058 103 2061 105
rect 2055 102 2061 103
rect 2065 137 2071 139
rect 2145 140 2150 142
rect 2145 138 2146 140
rect 2148 138 2150 140
rect 2065 135 2068 137
rect 2070 135 2071 137
rect 2065 134 2071 135
rect 2065 132 2068 134
rect 2070 132 2071 134
rect 2065 130 2071 132
rect 2065 128 2068 130
rect 2070 128 2071 130
rect 2065 126 2071 128
rect 2065 106 2069 126
rect 2081 129 2119 130
rect 2081 127 2116 129
rect 2118 127 2119 129
rect 2081 126 2119 127
rect 2114 123 2119 126
rect 2089 121 2104 122
rect 2089 119 2093 121
rect 2095 119 2100 121
rect 2102 119 2104 121
rect 2089 118 2104 119
rect 2114 121 2122 123
rect 2114 119 2119 121
rect 2121 119 2122 121
rect 2098 113 2102 118
rect 2114 117 2122 119
rect 2145 133 2150 138
rect 2145 131 2146 133
rect 2148 131 2150 133
rect 2145 129 2150 131
rect 2098 111 2099 113
rect 2101 111 2102 113
rect 2098 109 2102 111
rect 2065 105 2071 106
rect 2065 103 2068 105
rect 2070 103 2071 105
rect 2065 102 2071 103
rect 2146 111 2150 129
rect 2155 138 2159 139
rect 2155 136 2156 138
rect 2158 136 2159 138
rect 2155 130 2159 136
rect 2155 128 2176 130
rect 2155 126 2160 128
rect 2162 126 2176 128
rect 2146 109 2147 111
rect 2149 109 2150 111
rect 2155 121 2176 122
rect 2155 119 2156 121
rect 2158 119 2170 121
rect 2172 119 2176 121
rect 2155 118 2176 119
rect 2189 140 2191 142
rect 2187 135 2191 140
rect 2189 133 2191 135
rect 2199 141 2204 147
rect 2246 145 2259 146
rect 2246 143 2255 145
rect 2257 143 2259 145
rect 2199 139 2201 141
rect 2203 139 2204 141
rect 2246 142 2259 143
rect 2199 138 2204 139
rect 2199 134 2212 138
rect 2155 109 2159 118
rect 2187 117 2191 133
rect 2187 115 2188 117
rect 2190 115 2191 117
rect 2187 114 2191 115
rect 2186 112 2191 114
rect 2186 110 2187 112
rect 2189 110 2191 112
rect 2146 107 2150 109
rect 2186 108 2191 110
rect 2145 105 2150 107
rect 2145 103 2146 105
rect 2148 103 2150 105
rect 2213 121 2219 123
rect 2213 119 2214 121
rect 2216 119 2219 121
rect 2213 114 2219 119
rect 2206 113 2219 114
rect 2206 111 2207 113
rect 2209 111 2219 113
rect 2231 129 2243 131
rect 2231 127 2236 129
rect 2238 127 2243 129
rect 2231 126 2243 127
rect 2231 125 2241 126
rect 2239 124 2241 125
rect 2239 117 2243 124
rect 2206 110 2219 111
rect 2255 109 2259 142
rect 2267 141 2272 147
rect 2314 145 2327 146
rect 2314 143 2323 145
rect 2325 143 2327 145
rect 2267 139 2269 141
rect 2271 139 2272 141
rect 2314 142 2327 143
rect 2267 138 2272 139
rect 2267 134 2280 138
rect 2254 107 2259 109
rect 2145 101 2150 103
rect 2254 105 2255 107
rect 2257 105 2259 107
rect 2254 103 2259 105
rect 2281 121 2287 123
rect 2281 119 2282 121
rect 2284 119 2287 121
rect 2281 114 2287 119
rect 2274 113 2287 114
rect 2274 111 2276 113
rect 2278 111 2287 113
rect 2299 130 2311 131
rect 2299 128 2300 130
rect 2302 128 2311 130
rect 2299 126 2311 128
rect 2299 125 2309 126
rect 2307 124 2309 125
rect 2307 117 2311 124
rect 2274 110 2287 111
rect 2323 109 2327 142
rect 2322 107 2327 109
rect 2255 101 2259 103
rect 2322 105 2323 107
rect 2325 105 2327 107
rect 2322 103 2327 105
rect 2323 101 2327 103
rect 4 95 2331 96
rect 4 93 29 95
rect 31 93 39 95
rect 41 93 69 95
rect 71 93 79 95
rect 81 93 298 95
rect 300 93 336 95
rect 338 93 346 95
rect 348 93 565 95
rect 567 93 603 95
rect 605 93 613 95
rect 615 93 832 95
rect 834 93 870 95
rect 872 93 880 95
rect 882 93 1099 95
rect 1101 93 1137 95
rect 1139 93 1147 95
rect 1149 93 1366 95
rect 1368 93 1404 95
rect 1406 93 1414 95
rect 1416 93 1633 95
rect 1635 93 1671 95
rect 1673 93 1681 95
rect 1683 93 1900 95
rect 1902 93 1915 95
rect 1917 93 1968 95
rect 1970 93 2186 95
rect 2188 93 2331 95
rect 4 89 2331 93
rect 4 87 2276 89
rect 2278 87 2331 89
rect 4 85 2331 87
rect 4 83 2311 85
rect 2313 83 2331 85
rect 4 81 29 83
rect 31 81 39 83
rect 41 81 69 83
rect 71 81 79 83
rect 81 81 298 83
rect 300 81 336 83
rect 338 81 346 83
rect 348 81 565 83
rect 567 81 603 83
rect 605 81 613 83
rect 615 81 832 83
rect 834 81 870 83
rect 872 81 880 83
rect 882 81 1099 83
rect 1101 81 1137 83
rect 1139 81 1147 83
rect 1149 81 1366 83
rect 1368 81 1404 83
rect 1406 81 1414 83
rect 1416 81 1633 83
rect 1635 81 1671 83
rect 1673 81 1681 83
rect 1683 81 1900 83
rect 1902 81 1915 83
rect 1917 81 1968 83
rect 1970 81 2186 83
rect 2188 81 2331 83
rect 4 80 2331 81
rect 15 61 20 67
rect 32 71 44 75
rect 32 69 40 71
rect 42 69 44 71
rect 15 59 17 61
rect 19 59 20 61
rect 15 58 20 59
rect 15 57 29 58
rect 15 55 23 57
rect 25 55 29 57
rect 15 54 29 55
rect 8 49 21 50
rect 8 47 13 49
rect 15 47 21 49
rect 8 46 21 47
rect 8 37 12 46
rect 40 49 44 69
rect 55 58 60 67
rect 72 71 84 75
rect 72 69 80 71
rect 82 69 84 71
rect 55 57 69 58
rect 55 55 63 57
rect 65 55 69 57
rect 55 54 69 55
rect 39 47 41 49
rect 43 47 44 49
rect 39 44 44 47
rect 39 42 40 44
rect 42 42 44 44
rect 39 37 44 42
rect 48 49 61 50
rect 48 47 53 49
rect 55 47 61 49
rect 48 46 61 47
rect 48 41 52 46
rect 80 57 84 69
rect 80 55 81 57
rect 83 55 84 57
rect 80 49 84 55
rect 48 39 49 41
rect 51 39 52 41
rect 48 38 52 39
rect 79 47 84 49
rect 79 45 80 47
rect 82 45 84 47
rect 79 40 84 45
rect 39 35 40 37
rect 42 35 44 37
rect 39 33 44 35
rect 79 38 80 40
rect 82 38 84 40
rect 79 36 84 38
rect 88 73 93 75
rect 88 71 90 73
rect 92 71 93 73
rect 88 69 93 71
rect 88 65 92 69
rect 88 63 89 65
rect 91 63 92 65
rect 88 47 92 63
rect 167 73 173 74
rect 167 71 168 73
rect 170 71 173 73
rect 167 70 173 71
rect 88 45 93 47
rect 88 43 90 45
rect 92 43 93 45
rect 88 38 93 43
rect 116 57 124 59
rect 136 58 140 67
rect 116 55 117 57
rect 119 55 124 57
rect 116 53 124 55
rect 134 57 149 58
rect 134 55 136 57
rect 138 55 139 57
rect 141 55 143 57
rect 145 55 149 57
rect 134 54 149 55
rect 119 50 124 53
rect 169 57 173 70
rect 169 55 170 57
rect 172 55 173 57
rect 119 49 157 50
rect 119 47 133 49
rect 135 47 157 49
rect 119 46 157 47
rect 169 50 173 55
rect 167 48 173 50
rect 167 46 168 48
rect 170 46 173 48
rect 167 41 173 46
rect 167 39 168 41
rect 170 39 173 41
rect 88 36 90 38
rect 92 36 93 38
rect 88 34 93 36
rect 167 37 173 39
rect 177 73 183 74
rect 177 71 180 73
rect 182 71 183 73
rect 177 70 183 71
rect 257 74 264 75
rect 257 73 261 74
rect 257 71 258 73
rect 260 72 261 73
rect 263 72 264 74
rect 260 71 264 72
rect 177 50 181 70
rect 210 65 214 67
rect 210 63 211 65
rect 213 63 214 65
rect 177 48 183 50
rect 177 46 180 48
rect 182 46 183 48
rect 177 44 183 46
rect 177 42 180 44
rect 182 42 183 44
rect 177 41 183 42
rect 177 39 180 41
rect 182 39 183 41
rect 177 37 183 39
rect 210 58 214 63
rect 257 69 264 71
rect 201 57 216 58
rect 201 55 205 57
rect 207 55 212 57
rect 214 55 216 57
rect 201 54 216 55
rect 226 57 234 59
rect 226 55 231 57
rect 233 55 234 57
rect 226 53 234 55
rect 226 52 231 53
rect 226 50 228 52
rect 230 50 231 52
rect 193 46 231 50
rect 258 47 262 69
rect 267 63 271 64
rect 267 61 268 63
rect 270 61 271 63
rect 267 58 271 61
rect 267 57 288 58
rect 267 55 282 57
rect 284 55 288 57
rect 267 54 288 55
rect 298 66 303 68
rect 298 64 299 66
rect 301 64 303 66
rect 298 62 303 64
rect 257 45 262 47
rect 257 43 258 45
rect 260 43 262 45
rect 257 38 262 43
rect 257 36 258 38
rect 260 36 262 38
rect 267 48 272 50
rect 274 48 288 50
rect 267 46 288 48
rect 267 44 271 46
rect 267 42 268 44
rect 270 42 271 44
rect 267 37 271 42
rect 257 34 262 36
rect 299 43 303 62
rect 322 58 327 67
rect 339 71 351 75
rect 339 69 347 71
rect 349 69 351 71
rect 322 57 336 58
rect 322 55 330 57
rect 332 55 336 57
rect 322 54 336 55
rect 301 41 303 43
rect 299 36 303 41
rect 315 49 328 50
rect 315 47 320 49
rect 322 47 328 49
rect 315 46 328 47
rect 315 41 319 46
rect 347 57 351 69
rect 347 55 348 57
rect 350 55 351 57
rect 347 49 351 55
rect 315 39 316 41
rect 318 39 319 41
rect 315 38 319 39
rect 346 47 351 49
rect 346 45 347 47
rect 349 45 351 47
rect 346 40 351 45
rect 301 34 303 36
rect 290 33 303 34
rect 290 31 291 33
rect 293 31 303 33
rect 290 30 303 31
rect 299 29 303 30
rect 346 38 347 40
rect 349 38 351 40
rect 346 36 351 38
rect 355 73 360 75
rect 355 71 357 73
rect 359 71 360 73
rect 355 69 360 71
rect 355 65 359 69
rect 355 63 356 65
rect 358 63 359 65
rect 355 47 359 63
rect 434 73 440 74
rect 434 71 435 73
rect 437 71 440 73
rect 434 70 440 71
rect 355 45 360 47
rect 355 43 357 45
rect 359 43 360 45
rect 355 38 360 43
rect 383 57 391 59
rect 403 58 407 67
rect 383 55 384 57
rect 386 55 391 57
rect 383 53 391 55
rect 401 57 416 58
rect 401 55 403 57
rect 405 55 406 57
rect 408 55 410 57
rect 412 55 416 57
rect 401 54 416 55
rect 386 50 391 53
rect 436 57 440 70
rect 436 55 437 57
rect 439 55 440 57
rect 386 49 424 50
rect 386 47 400 49
rect 402 47 424 49
rect 386 46 424 47
rect 436 50 440 55
rect 434 48 440 50
rect 434 46 435 48
rect 437 46 440 48
rect 434 41 440 46
rect 434 39 435 41
rect 437 39 440 41
rect 355 36 357 38
rect 359 36 360 38
rect 355 34 360 36
rect 434 37 440 39
rect 444 73 450 74
rect 444 71 447 73
rect 449 71 450 73
rect 444 70 450 71
rect 524 74 531 75
rect 524 73 528 74
rect 524 71 525 73
rect 527 72 528 73
rect 530 72 531 74
rect 527 71 531 72
rect 444 50 448 70
rect 477 65 481 67
rect 477 63 478 65
rect 480 63 481 65
rect 444 48 450 50
rect 444 46 447 48
rect 449 46 450 48
rect 444 44 450 46
rect 444 42 447 44
rect 449 42 450 44
rect 444 41 450 42
rect 444 39 447 41
rect 449 39 450 41
rect 444 37 450 39
rect 477 58 481 63
rect 524 69 531 71
rect 468 57 483 58
rect 468 55 472 57
rect 474 55 479 57
rect 481 55 483 57
rect 468 54 483 55
rect 493 57 501 59
rect 493 55 498 57
rect 500 55 501 57
rect 493 53 501 55
rect 493 52 498 53
rect 493 50 495 52
rect 497 50 498 52
rect 460 46 498 50
rect 525 47 529 69
rect 534 63 538 64
rect 534 61 535 63
rect 537 61 538 63
rect 534 58 538 61
rect 534 57 555 58
rect 534 55 549 57
rect 551 55 555 57
rect 534 54 555 55
rect 565 66 570 68
rect 565 64 566 66
rect 568 64 570 66
rect 565 62 570 64
rect 524 45 529 47
rect 524 43 525 45
rect 527 43 529 45
rect 524 38 529 43
rect 524 36 525 38
rect 527 36 529 38
rect 534 48 539 50
rect 541 48 555 50
rect 534 46 555 48
rect 534 44 538 46
rect 534 42 535 44
rect 537 42 538 44
rect 534 37 538 42
rect 524 34 529 36
rect 566 43 570 62
rect 589 58 594 67
rect 606 71 618 75
rect 606 69 614 71
rect 616 69 618 71
rect 589 57 603 58
rect 589 55 597 57
rect 599 55 603 57
rect 589 54 603 55
rect 568 41 570 43
rect 566 36 570 41
rect 582 49 595 50
rect 582 47 587 49
rect 589 47 595 49
rect 582 46 595 47
rect 582 41 586 46
rect 614 57 618 69
rect 614 55 615 57
rect 617 55 618 57
rect 614 49 618 55
rect 582 39 583 41
rect 585 39 586 41
rect 582 38 586 39
rect 613 47 618 49
rect 613 45 614 47
rect 616 45 618 47
rect 613 40 618 45
rect 568 34 570 36
rect 557 33 570 34
rect 557 31 558 33
rect 560 31 570 33
rect 557 30 570 31
rect 566 29 570 30
rect 613 38 614 40
rect 616 38 618 40
rect 613 36 618 38
rect 622 73 627 75
rect 622 71 624 73
rect 626 71 627 73
rect 622 69 627 71
rect 622 65 626 69
rect 622 63 623 65
rect 625 63 626 65
rect 622 47 626 63
rect 701 73 707 74
rect 701 71 702 73
rect 704 71 707 73
rect 701 70 707 71
rect 622 45 627 47
rect 622 43 624 45
rect 626 43 627 45
rect 622 38 627 43
rect 650 57 658 59
rect 670 58 674 67
rect 650 55 651 57
rect 653 55 658 57
rect 650 53 658 55
rect 668 57 683 58
rect 668 55 670 57
rect 672 55 673 57
rect 675 55 677 57
rect 679 55 683 57
rect 668 54 683 55
rect 653 50 658 53
rect 703 57 707 70
rect 703 55 704 57
rect 706 55 707 57
rect 653 49 691 50
rect 653 47 667 49
rect 669 47 691 49
rect 653 46 691 47
rect 703 50 707 55
rect 701 48 707 50
rect 701 46 702 48
rect 704 46 707 48
rect 701 41 707 46
rect 701 39 702 41
rect 704 39 707 41
rect 622 36 624 38
rect 626 36 627 38
rect 622 34 627 36
rect 701 37 707 39
rect 711 73 717 74
rect 711 71 714 73
rect 716 71 717 73
rect 711 70 717 71
rect 791 74 798 75
rect 791 73 795 74
rect 791 71 792 73
rect 794 72 795 73
rect 797 72 798 74
rect 794 71 798 72
rect 711 50 715 70
rect 744 65 748 67
rect 744 63 745 65
rect 747 63 748 65
rect 711 48 717 50
rect 711 46 714 48
rect 716 46 717 48
rect 711 44 717 46
rect 711 42 714 44
rect 716 42 717 44
rect 711 41 717 42
rect 711 39 714 41
rect 716 39 717 41
rect 711 37 717 39
rect 744 58 748 63
rect 791 69 798 71
rect 735 57 750 58
rect 735 55 739 57
rect 741 55 746 57
rect 748 55 750 57
rect 735 54 750 55
rect 760 57 768 59
rect 760 55 765 57
rect 767 55 768 57
rect 760 53 768 55
rect 760 52 765 53
rect 760 50 762 52
rect 764 50 765 52
rect 727 46 765 50
rect 792 47 796 69
rect 801 63 805 64
rect 801 61 802 63
rect 804 61 805 63
rect 801 58 805 61
rect 801 57 822 58
rect 801 55 816 57
rect 818 55 822 57
rect 801 54 822 55
rect 832 66 837 68
rect 832 64 833 66
rect 835 64 837 66
rect 832 62 837 64
rect 791 45 796 47
rect 791 43 792 45
rect 794 43 796 45
rect 791 38 796 43
rect 791 36 792 38
rect 794 36 796 38
rect 801 48 806 50
rect 808 48 822 50
rect 801 46 822 48
rect 801 44 805 46
rect 801 42 802 44
rect 804 42 805 44
rect 801 37 805 42
rect 791 34 796 36
rect 833 43 837 62
rect 856 58 861 67
rect 873 71 885 75
rect 873 69 881 71
rect 883 69 885 71
rect 856 57 870 58
rect 856 55 864 57
rect 866 55 870 57
rect 856 54 870 55
rect 835 41 837 43
rect 833 36 837 41
rect 849 49 862 50
rect 849 47 854 49
rect 856 47 862 49
rect 849 46 862 47
rect 849 41 853 46
rect 881 57 885 69
rect 881 55 882 57
rect 884 55 885 57
rect 881 49 885 55
rect 849 39 850 41
rect 852 39 853 41
rect 849 38 853 39
rect 880 47 885 49
rect 880 45 881 47
rect 883 45 885 47
rect 880 40 885 45
rect 835 34 837 36
rect 824 33 837 34
rect 824 31 825 33
rect 827 31 837 33
rect 824 30 837 31
rect 833 29 837 30
rect 880 38 881 40
rect 883 38 885 40
rect 880 36 885 38
rect 889 73 894 75
rect 889 71 891 73
rect 893 71 894 73
rect 889 69 894 71
rect 889 65 893 69
rect 889 63 890 65
rect 892 63 893 65
rect 889 47 893 63
rect 968 73 974 74
rect 968 71 969 73
rect 971 71 974 73
rect 968 70 974 71
rect 889 45 894 47
rect 889 43 891 45
rect 893 43 894 45
rect 889 38 894 43
rect 917 57 925 59
rect 937 58 941 67
rect 917 55 918 57
rect 920 55 925 57
rect 917 53 925 55
rect 935 57 950 58
rect 935 55 937 57
rect 939 55 940 57
rect 942 55 944 57
rect 946 55 950 57
rect 935 54 950 55
rect 920 50 925 53
rect 970 57 974 70
rect 970 55 971 57
rect 973 55 974 57
rect 920 49 958 50
rect 920 47 934 49
rect 936 47 958 49
rect 920 46 958 47
rect 970 50 974 55
rect 968 48 974 50
rect 968 46 969 48
rect 971 46 974 48
rect 968 41 974 46
rect 968 39 969 41
rect 971 39 974 41
rect 889 36 891 38
rect 893 36 894 38
rect 889 34 894 36
rect 968 37 974 39
rect 978 73 984 74
rect 978 71 981 73
rect 983 71 984 73
rect 978 70 984 71
rect 1058 74 1065 75
rect 1058 73 1062 74
rect 1058 71 1059 73
rect 1061 72 1062 73
rect 1064 72 1065 74
rect 1061 71 1065 72
rect 978 50 982 70
rect 1011 65 1015 67
rect 1011 63 1012 65
rect 1014 63 1015 65
rect 978 48 984 50
rect 978 46 981 48
rect 983 46 984 48
rect 978 44 984 46
rect 978 42 981 44
rect 983 42 984 44
rect 978 41 984 42
rect 978 39 981 41
rect 983 39 984 41
rect 978 37 984 39
rect 1011 58 1015 63
rect 1058 69 1065 71
rect 1002 57 1017 58
rect 1002 55 1006 57
rect 1008 55 1013 57
rect 1015 55 1017 57
rect 1002 54 1017 55
rect 1027 57 1035 59
rect 1027 55 1032 57
rect 1034 55 1035 57
rect 1027 53 1035 55
rect 1027 52 1032 53
rect 1027 50 1029 52
rect 1031 50 1032 52
rect 994 46 1032 50
rect 1059 47 1063 69
rect 1068 63 1072 64
rect 1068 61 1069 63
rect 1071 61 1072 63
rect 1068 58 1072 61
rect 1068 57 1089 58
rect 1068 55 1083 57
rect 1085 55 1089 57
rect 1068 54 1089 55
rect 1099 66 1104 68
rect 1099 64 1100 66
rect 1102 64 1104 66
rect 1099 62 1104 64
rect 1058 45 1063 47
rect 1058 43 1059 45
rect 1061 43 1063 45
rect 1058 38 1063 43
rect 1058 36 1059 38
rect 1061 36 1063 38
rect 1068 48 1073 50
rect 1075 48 1089 50
rect 1068 46 1089 48
rect 1068 44 1072 46
rect 1068 42 1069 44
rect 1071 42 1072 44
rect 1068 37 1072 42
rect 1058 34 1063 36
rect 1100 43 1104 62
rect 1123 58 1128 67
rect 1140 71 1152 75
rect 1140 69 1148 71
rect 1150 69 1152 71
rect 1123 57 1137 58
rect 1123 55 1131 57
rect 1133 55 1137 57
rect 1123 54 1137 55
rect 1102 41 1104 43
rect 1100 36 1104 41
rect 1116 49 1129 50
rect 1116 47 1121 49
rect 1123 47 1129 49
rect 1116 46 1129 47
rect 1116 41 1120 46
rect 1148 57 1152 69
rect 1148 55 1149 57
rect 1151 55 1152 57
rect 1148 49 1152 55
rect 1116 39 1117 41
rect 1119 39 1120 41
rect 1116 38 1120 39
rect 1147 47 1152 49
rect 1147 45 1148 47
rect 1150 45 1152 47
rect 1147 40 1152 45
rect 1102 34 1104 36
rect 1091 33 1104 34
rect 1091 31 1092 33
rect 1094 31 1104 33
rect 1091 30 1104 31
rect 1100 29 1104 30
rect 1147 38 1148 40
rect 1150 38 1152 40
rect 1147 36 1152 38
rect 1156 73 1161 75
rect 1156 71 1158 73
rect 1160 71 1161 73
rect 1156 69 1161 71
rect 1156 65 1160 69
rect 1156 63 1157 65
rect 1159 63 1160 65
rect 1156 47 1160 63
rect 1235 73 1241 74
rect 1235 71 1236 73
rect 1238 71 1241 73
rect 1235 70 1241 71
rect 1156 45 1161 47
rect 1156 43 1158 45
rect 1160 43 1161 45
rect 1156 38 1161 43
rect 1184 57 1192 59
rect 1204 58 1208 67
rect 1184 55 1185 57
rect 1187 55 1192 57
rect 1184 53 1192 55
rect 1202 57 1217 58
rect 1202 55 1204 57
rect 1206 55 1207 57
rect 1209 55 1211 57
rect 1213 55 1217 57
rect 1202 54 1217 55
rect 1187 50 1192 53
rect 1237 57 1241 70
rect 1237 55 1238 57
rect 1240 55 1241 57
rect 1187 49 1225 50
rect 1187 47 1201 49
rect 1203 47 1225 49
rect 1187 46 1225 47
rect 1237 50 1241 55
rect 1235 48 1241 50
rect 1235 46 1236 48
rect 1238 46 1241 48
rect 1235 41 1241 46
rect 1235 39 1236 41
rect 1238 39 1241 41
rect 1156 36 1158 38
rect 1160 36 1161 38
rect 1156 34 1161 36
rect 1235 37 1241 39
rect 1245 73 1251 74
rect 1245 71 1248 73
rect 1250 71 1251 73
rect 1245 70 1251 71
rect 1325 74 1332 75
rect 1325 73 1329 74
rect 1325 71 1326 73
rect 1328 72 1329 73
rect 1331 72 1332 74
rect 1328 71 1332 72
rect 1245 50 1249 70
rect 1278 65 1282 67
rect 1278 63 1279 65
rect 1281 63 1282 65
rect 1245 48 1251 50
rect 1245 46 1248 48
rect 1250 46 1251 48
rect 1245 44 1251 46
rect 1245 42 1248 44
rect 1250 42 1251 44
rect 1245 41 1251 42
rect 1245 39 1248 41
rect 1250 39 1251 41
rect 1245 37 1251 39
rect 1278 58 1282 63
rect 1325 69 1332 71
rect 1269 57 1284 58
rect 1269 55 1273 57
rect 1275 55 1280 57
rect 1282 55 1284 57
rect 1269 54 1284 55
rect 1294 57 1302 59
rect 1294 55 1299 57
rect 1301 55 1302 57
rect 1294 53 1302 55
rect 1294 52 1299 53
rect 1294 50 1296 52
rect 1298 50 1299 52
rect 1261 46 1299 50
rect 1326 47 1330 69
rect 1335 63 1339 64
rect 1335 61 1336 63
rect 1338 61 1339 63
rect 1335 58 1339 61
rect 1335 57 1356 58
rect 1335 55 1350 57
rect 1352 55 1356 57
rect 1335 54 1356 55
rect 1366 66 1371 68
rect 1366 64 1367 66
rect 1369 64 1371 66
rect 1366 62 1371 64
rect 1325 45 1330 47
rect 1325 43 1326 45
rect 1328 43 1330 45
rect 1325 38 1330 43
rect 1325 36 1326 38
rect 1328 36 1330 38
rect 1335 48 1340 50
rect 1342 48 1356 50
rect 1335 46 1356 48
rect 1335 44 1339 46
rect 1335 42 1336 44
rect 1338 42 1339 44
rect 1335 37 1339 42
rect 1325 34 1330 36
rect 1367 43 1371 62
rect 1390 58 1395 67
rect 1407 71 1419 75
rect 1407 69 1415 71
rect 1417 69 1419 71
rect 1390 57 1404 58
rect 1390 55 1398 57
rect 1400 55 1404 57
rect 1390 54 1404 55
rect 1369 41 1371 43
rect 1367 36 1371 41
rect 1383 49 1396 50
rect 1383 47 1388 49
rect 1390 47 1396 49
rect 1383 46 1396 47
rect 1383 41 1387 46
rect 1415 57 1419 69
rect 1415 55 1416 57
rect 1418 55 1419 57
rect 1415 49 1419 55
rect 1383 39 1384 41
rect 1386 39 1387 41
rect 1383 38 1387 39
rect 1414 47 1419 49
rect 1414 45 1415 47
rect 1417 45 1419 47
rect 1414 40 1419 45
rect 1369 34 1371 36
rect 1358 33 1371 34
rect 1358 31 1359 33
rect 1361 31 1371 33
rect 1358 30 1371 31
rect 1367 29 1371 30
rect 1414 38 1415 40
rect 1417 38 1419 40
rect 1414 36 1419 38
rect 1423 73 1428 75
rect 1423 71 1425 73
rect 1427 71 1428 73
rect 1423 69 1428 71
rect 1423 65 1427 69
rect 1423 63 1424 65
rect 1426 63 1427 65
rect 1423 47 1427 63
rect 1502 73 1508 74
rect 1502 71 1503 73
rect 1505 71 1508 73
rect 1502 70 1508 71
rect 1423 45 1428 47
rect 1423 43 1425 45
rect 1427 43 1428 45
rect 1423 38 1428 43
rect 1451 57 1459 59
rect 1471 58 1475 67
rect 1451 55 1452 57
rect 1454 55 1459 57
rect 1451 53 1459 55
rect 1469 57 1484 58
rect 1469 55 1471 57
rect 1473 55 1474 57
rect 1476 55 1478 57
rect 1480 55 1484 57
rect 1469 54 1484 55
rect 1454 50 1459 53
rect 1504 57 1508 70
rect 1504 55 1505 57
rect 1507 55 1508 57
rect 1454 49 1492 50
rect 1454 47 1468 49
rect 1470 47 1492 49
rect 1454 46 1492 47
rect 1504 50 1508 55
rect 1502 48 1508 50
rect 1502 46 1503 48
rect 1505 46 1508 48
rect 1502 41 1508 46
rect 1502 39 1503 41
rect 1505 39 1508 41
rect 1423 36 1425 38
rect 1427 36 1428 38
rect 1423 34 1428 36
rect 1502 37 1508 39
rect 1512 73 1518 74
rect 1512 71 1515 73
rect 1517 71 1518 73
rect 1512 70 1518 71
rect 1592 74 1599 75
rect 1592 73 1596 74
rect 1592 71 1593 73
rect 1595 72 1596 73
rect 1598 72 1599 74
rect 1595 71 1599 72
rect 1512 50 1516 70
rect 1545 65 1549 67
rect 1545 63 1546 65
rect 1548 63 1549 65
rect 1512 48 1518 50
rect 1512 46 1515 48
rect 1517 46 1518 48
rect 1512 44 1518 46
rect 1512 42 1515 44
rect 1517 42 1518 44
rect 1512 41 1518 42
rect 1512 39 1515 41
rect 1517 39 1518 41
rect 1512 37 1518 39
rect 1545 58 1549 63
rect 1592 69 1599 71
rect 1536 57 1551 58
rect 1536 55 1540 57
rect 1542 55 1547 57
rect 1549 55 1551 57
rect 1536 54 1551 55
rect 1561 57 1569 59
rect 1561 55 1566 57
rect 1568 55 1569 57
rect 1561 53 1569 55
rect 1561 52 1566 53
rect 1561 50 1563 52
rect 1565 50 1566 52
rect 1528 46 1566 50
rect 1593 47 1597 69
rect 1602 63 1606 64
rect 1602 61 1603 63
rect 1605 61 1606 63
rect 1602 58 1606 61
rect 1602 57 1623 58
rect 1602 55 1617 57
rect 1619 55 1623 57
rect 1602 54 1623 55
rect 1633 66 1638 68
rect 1633 64 1634 66
rect 1636 64 1638 66
rect 1633 62 1638 64
rect 1592 45 1597 47
rect 1592 43 1593 45
rect 1595 43 1597 45
rect 1592 38 1597 43
rect 1592 36 1593 38
rect 1595 36 1597 38
rect 1602 48 1607 50
rect 1609 48 1623 50
rect 1602 46 1623 48
rect 1602 44 1606 46
rect 1602 42 1603 44
rect 1605 42 1606 44
rect 1602 37 1606 42
rect 1592 34 1597 36
rect 1634 43 1638 62
rect 1657 58 1662 67
rect 1674 71 1686 75
rect 1674 69 1682 71
rect 1684 69 1686 71
rect 1657 57 1671 58
rect 1657 55 1665 57
rect 1667 55 1671 57
rect 1657 54 1671 55
rect 1636 41 1638 43
rect 1634 36 1638 41
rect 1650 49 1663 50
rect 1650 47 1655 49
rect 1657 47 1663 49
rect 1650 46 1663 47
rect 1650 41 1654 46
rect 1682 57 1686 69
rect 1682 55 1683 57
rect 1685 55 1686 57
rect 1682 49 1686 55
rect 1650 39 1651 41
rect 1653 39 1654 41
rect 1650 38 1654 39
rect 1681 47 1686 49
rect 1681 45 1682 47
rect 1684 45 1686 47
rect 1681 40 1686 45
rect 1636 34 1638 36
rect 1625 33 1638 34
rect 1625 31 1626 33
rect 1628 31 1638 33
rect 1625 30 1638 31
rect 1634 29 1638 30
rect 1681 38 1682 40
rect 1684 38 1686 40
rect 1681 36 1686 38
rect 1690 73 1695 75
rect 1690 71 1692 73
rect 1694 71 1695 73
rect 1690 69 1695 71
rect 1690 65 1694 69
rect 1690 63 1691 65
rect 1693 63 1694 65
rect 1690 47 1694 63
rect 1769 73 1775 74
rect 1769 71 1770 73
rect 1772 71 1775 73
rect 1769 70 1775 71
rect 1690 45 1695 47
rect 1690 43 1692 45
rect 1694 43 1695 45
rect 1690 38 1695 43
rect 1718 57 1726 59
rect 1738 58 1742 67
rect 1718 55 1719 57
rect 1721 55 1726 57
rect 1718 53 1726 55
rect 1736 57 1751 58
rect 1736 55 1738 57
rect 1740 55 1741 57
rect 1743 55 1745 57
rect 1747 55 1751 57
rect 1736 54 1751 55
rect 1721 50 1726 53
rect 1771 57 1775 70
rect 1771 55 1772 57
rect 1774 55 1775 57
rect 1721 49 1759 50
rect 1721 47 1735 49
rect 1737 47 1759 49
rect 1721 46 1759 47
rect 1771 50 1775 55
rect 1769 48 1775 50
rect 1769 46 1770 48
rect 1772 46 1775 48
rect 1769 41 1775 46
rect 1769 39 1770 41
rect 1772 39 1775 41
rect 1690 36 1692 38
rect 1694 36 1695 38
rect 1690 34 1695 36
rect 1769 37 1775 39
rect 1779 73 1785 74
rect 1779 71 1782 73
rect 1784 71 1785 73
rect 1779 70 1785 71
rect 1859 74 1866 75
rect 1859 73 1863 74
rect 1859 71 1860 73
rect 1862 72 1863 73
rect 1865 72 1866 74
rect 1862 71 1866 72
rect 1948 73 1972 74
rect 1779 50 1783 70
rect 1812 65 1816 67
rect 1812 63 1813 65
rect 1815 63 1816 65
rect 1779 48 1785 50
rect 1779 46 1782 48
rect 1784 46 1785 48
rect 1779 44 1785 46
rect 1779 42 1782 44
rect 1784 42 1785 44
rect 1779 41 1785 42
rect 1779 39 1782 41
rect 1784 39 1785 41
rect 1779 37 1785 39
rect 1812 58 1816 63
rect 1859 69 1866 71
rect 1948 71 1950 73
rect 1952 71 1972 73
rect 1948 70 1972 71
rect 1803 57 1818 58
rect 1803 55 1807 57
rect 1809 55 1814 57
rect 1816 55 1818 57
rect 1803 54 1818 55
rect 1828 57 1836 59
rect 1828 55 1833 57
rect 1835 55 1836 57
rect 1828 53 1836 55
rect 1828 52 1833 53
rect 1828 50 1830 52
rect 1832 50 1833 52
rect 1795 46 1833 50
rect 1860 47 1864 69
rect 1869 63 1873 64
rect 1869 61 1870 63
rect 1872 61 1873 63
rect 1869 58 1873 61
rect 1869 57 1890 58
rect 1869 55 1884 57
rect 1886 55 1890 57
rect 1869 54 1890 55
rect 1900 66 1905 68
rect 1900 64 1901 66
rect 1903 64 1905 66
rect 1900 62 1905 64
rect 1859 45 1864 47
rect 1859 43 1860 45
rect 1862 43 1864 45
rect 1859 38 1864 43
rect 1859 36 1860 38
rect 1862 36 1864 38
rect 1869 48 1874 50
rect 1876 48 1890 50
rect 1869 46 1890 48
rect 1869 44 1873 46
rect 1869 42 1870 44
rect 1872 42 1873 44
rect 1869 37 1873 42
rect 1859 34 1864 36
rect 1901 43 1905 62
rect 1920 66 1933 67
rect 1920 64 1925 66
rect 1927 64 1933 66
rect 1920 62 1933 64
rect 1920 61 1930 62
rect 1928 60 1930 61
rect 1932 60 1933 62
rect 1903 41 1905 43
rect 1901 36 1905 41
rect 1903 34 1905 36
rect 1892 33 1905 34
rect 1892 31 1893 33
rect 1895 31 1905 33
rect 1892 30 1905 31
rect 1901 29 1905 30
rect 1912 49 1917 51
rect 1912 47 1914 49
rect 1916 47 1917 49
rect 1912 35 1917 47
rect 1928 53 1933 60
rect 1912 29 1924 35
rect 1968 49 1972 70
rect 1968 47 1969 49
rect 1971 47 1972 49
rect 1968 42 1972 47
rect 1956 40 1972 42
rect 1956 38 1958 40
rect 1960 38 1972 40
rect 1956 37 1972 38
rect 1976 73 1981 75
rect 1976 71 1978 73
rect 1980 71 1981 73
rect 1976 69 1981 71
rect 1976 65 1980 69
rect 1976 63 1977 65
rect 1979 63 1980 65
rect 1976 47 1980 63
rect 2055 73 2061 74
rect 2055 71 2056 73
rect 2058 71 2061 73
rect 2055 70 2061 71
rect 1976 45 1981 47
rect 1976 43 1978 45
rect 1980 43 1981 45
rect 1976 38 1981 43
rect 2004 57 2012 59
rect 2024 58 2028 67
rect 2004 55 2005 57
rect 2007 55 2012 57
rect 2004 53 2012 55
rect 2022 57 2037 58
rect 2022 55 2024 57
rect 2026 55 2031 57
rect 2033 55 2037 57
rect 2022 54 2037 55
rect 2007 50 2012 53
rect 2057 57 2061 70
rect 2057 55 2058 57
rect 2060 55 2061 57
rect 2007 49 2045 50
rect 2007 47 2018 49
rect 2020 47 2045 49
rect 2007 46 2045 47
rect 2057 50 2061 55
rect 2055 48 2061 50
rect 2055 46 2056 48
rect 2058 46 2061 48
rect 2055 41 2061 46
rect 2055 39 2056 41
rect 2058 39 2061 41
rect 1976 36 1978 38
rect 1980 36 1981 38
rect 1976 34 1981 36
rect 2055 37 2061 39
rect 2065 73 2071 74
rect 2065 71 2068 73
rect 2070 71 2071 73
rect 2065 70 2071 71
rect 2145 74 2152 75
rect 2145 73 2149 74
rect 2145 71 2146 73
rect 2148 72 2149 73
rect 2151 72 2152 74
rect 2148 71 2152 72
rect 2065 50 2069 70
rect 2098 65 2102 67
rect 2098 63 2099 65
rect 2101 63 2102 65
rect 2065 48 2071 50
rect 2065 46 2068 48
rect 2070 46 2071 48
rect 2065 44 2071 46
rect 2065 42 2068 44
rect 2070 42 2071 44
rect 2065 41 2071 42
rect 2065 39 2068 41
rect 2070 39 2071 41
rect 2065 37 2071 39
rect 2098 58 2102 63
rect 2145 69 2151 71
rect 2089 57 2104 58
rect 2089 55 2093 57
rect 2095 55 2100 57
rect 2102 55 2104 57
rect 2089 54 2104 55
rect 2114 57 2122 59
rect 2114 55 2119 57
rect 2121 55 2122 57
rect 2114 53 2122 55
rect 2114 52 2119 53
rect 2114 50 2116 52
rect 2118 50 2119 52
rect 2081 46 2119 50
rect 2146 47 2150 69
rect 2155 63 2159 67
rect 2155 61 2156 63
rect 2158 61 2159 63
rect 2155 58 2159 61
rect 2155 57 2176 58
rect 2155 55 2170 57
rect 2172 55 2176 57
rect 2155 54 2176 55
rect 2186 66 2191 68
rect 2186 64 2187 66
rect 2189 64 2191 66
rect 2186 62 2191 64
rect 2145 45 2150 47
rect 2145 43 2146 45
rect 2148 43 2150 45
rect 2145 38 2150 43
rect 2145 36 2146 38
rect 2148 36 2150 38
rect 2155 48 2160 50
rect 2162 48 2176 50
rect 2155 46 2176 48
rect 2155 44 2159 46
rect 2155 42 2156 44
rect 2158 42 2159 44
rect 2155 37 2159 42
rect 2145 34 2150 36
rect 2187 43 2191 62
rect 2255 73 2259 75
rect 2254 71 2259 73
rect 2254 69 2255 71
rect 2257 69 2259 71
rect 2254 67 2259 69
rect 2206 65 2219 66
rect 2206 63 2210 65
rect 2212 63 2219 65
rect 2206 62 2219 63
rect 2213 57 2219 62
rect 2213 55 2214 57
rect 2216 55 2219 57
rect 2213 53 2219 55
rect 2239 52 2243 59
rect 2239 51 2241 52
rect 2231 50 2241 51
rect 2231 48 2236 50
rect 2238 48 2243 50
rect 2231 45 2243 48
rect 2189 41 2191 43
rect 2187 36 2191 41
rect 2189 34 2191 36
rect 2178 33 2191 34
rect 2178 31 2180 33
rect 2182 31 2191 33
rect 2178 30 2191 31
rect 2187 29 2191 30
rect 2199 38 2212 42
rect 2199 37 2204 38
rect 2199 35 2201 37
rect 2203 35 2204 37
rect 2199 29 2204 35
rect 2255 34 2259 67
rect 2323 73 2327 75
rect 2322 71 2327 73
rect 2322 69 2323 71
rect 2325 69 2327 71
rect 2322 67 2327 69
rect 2274 65 2287 66
rect 2274 63 2276 65
rect 2278 63 2287 65
rect 2274 62 2287 63
rect 2281 57 2287 62
rect 2281 55 2282 57
rect 2284 55 2287 57
rect 2281 53 2287 55
rect 2307 52 2311 59
rect 2307 51 2309 52
rect 2299 50 2309 51
rect 2299 48 2300 50
rect 2302 48 2311 50
rect 2299 45 2311 48
rect 2246 33 2259 34
rect 2246 31 2255 33
rect 2257 31 2259 33
rect 2246 30 2259 31
rect 2267 38 2280 42
rect 2267 37 2272 38
rect 2267 35 2269 37
rect 2271 35 2272 37
rect 2267 29 2272 35
rect 2323 34 2327 67
rect 2314 33 2327 34
rect 2314 31 2323 33
rect 2325 31 2327 33
rect 2314 30 2327 31
rect 4 23 2331 24
rect 4 21 39 23
rect 41 21 79 23
rect 81 21 298 23
rect 300 21 346 23
rect 348 21 565 23
rect 567 21 613 23
rect 615 21 832 23
rect 834 21 880 23
rect 882 21 1099 23
rect 1101 21 1147 23
rect 1149 21 1366 23
rect 1368 21 1414 23
rect 1416 21 1633 23
rect 1635 21 1681 23
rect 1683 21 1900 23
rect 1902 21 1948 23
rect 1950 21 2186 23
rect 2188 21 2320 23
rect 2322 21 2331 23
rect 4 11 2331 21
rect 4 9 39 11
rect 41 9 79 11
rect 81 9 298 11
rect 300 9 346 11
rect 348 9 565 11
rect 567 9 613 11
rect 615 9 832 11
rect 834 9 880 11
rect 882 9 1099 11
rect 1101 9 1147 11
rect 1149 9 1366 11
rect 1368 9 1414 11
rect 1416 9 1633 11
rect 1635 9 1681 11
rect 1683 9 1900 11
rect 1902 9 1948 11
rect 1950 9 2186 11
rect 2188 9 2331 11
rect 4 8 2331 9
rect 8 -12 12 -5
rect 39 -6 44 -4
rect 8 -14 9 -12
rect 11 -14 12 -12
rect 8 -15 21 -14
rect 8 -17 13 -15
rect 15 -17 21 -15
rect 8 -18 21 -17
rect 15 -23 29 -22
rect 15 -25 23 -23
rect 25 -25 29 -23
rect 15 -26 29 -25
rect 39 -8 40 -6
rect 42 -8 44 -6
rect 39 -13 44 -8
rect 39 -15 40 -13
rect 42 -15 44 -13
rect 39 -17 44 -15
rect 15 -35 20 -26
rect 40 -18 44 -17
rect 48 -14 52 -5
rect 299 2 303 3
rect 290 -2 303 2
rect 88 -4 93 -2
rect 79 -6 84 -4
rect 48 -15 61 -14
rect 48 -17 53 -15
rect 55 -17 61 -15
rect 48 -18 61 -17
rect 40 -20 41 -18
rect 43 -20 44 -18
rect 40 -37 44 -20
rect 55 -23 69 -22
rect 55 -25 63 -23
rect 65 -25 69 -23
rect 55 -26 69 -25
rect 79 -8 80 -6
rect 82 -8 84 -6
rect 79 -13 84 -8
rect 79 -15 80 -13
rect 82 -15 84 -13
rect 79 -17 84 -15
rect 55 -29 60 -26
rect 55 -31 57 -29
rect 59 -31 60 -29
rect 55 -35 60 -31
rect 80 -23 84 -17
rect 80 -25 81 -23
rect 83 -25 84 -23
rect 32 -39 40 -37
rect 42 -39 44 -37
rect 80 -37 84 -25
rect 32 -43 44 -39
rect 72 -39 80 -37
rect 82 -39 84 -37
rect 72 -43 84 -39
rect 88 -6 90 -4
rect 92 -6 93 -4
rect 88 -11 93 -6
rect 88 -13 90 -11
rect 92 -13 93 -11
rect 88 -15 93 -13
rect 88 -31 92 -15
rect 119 -15 157 -14
rect 119 -17 121 -15
rect 123 -17 157 -15
rect 119 -18 157 -17
rect 119 -21 124 -18
rect 116 -23 124 -21
rect 116 -25 117 -23
rect 119 -25 124 -23
rect 116 -27 124 -25
rect 134 -23 149 -22
rect 134 -25 136 -23
rect 138 -25 139 -23
rect 141 -25 143 -23
rect 145 -25 149 -23
rect 134 -26 149 -25
rect 88 -33 89 -31
rect 91 -33 92 -31
rect 88 -37 92 -33
rect 88 -39 93 -37
rect 136 -35 140 -26
rect 167 -7 173 -5
rect 167 -9 168 -7
rect 170 -9 173 -7
rect 167 -14 173 -9
rect 167 -16 168 -14
rect 170 -16 173 -14
rect 167 -18 173 -16
rect 169 -23 173 -18
rect 169 -25 170 -23
rect 172 -25 173 -23
rect 169 -38 173 -25
rect 88 -41 90 -39
rect 92 -41 93 -39
rect 88 -43 93 -41
rect 167 -39 173 -38
rect 167 -41 168 -39
rect 170 -41 173 -39
rect 167 -42 173 -41
rect 177 -7 183 -5
rect 257 -4 262 -2
rect 257 -6 258 -4
rect 260 -6 262 -4
rect 177 -9 180 -7
rect 182 -9 183 -7
rect 177 -10 183 -9
rect 177 -12 180 -10
rect 182 -12 183 -10
rect 177 -14 183 -12
rect 177 -16 180 -14
rect 182 -16 183 -14
rect 177 -18 183 -16
rect 177 -38 181 -18
rect 193 -15 231 -14
rect 193 -17 227 -15
rect 229 -17 231 -15
rect 193 -18 231 -17
rect 226 -21 231 -18
rect 201 -23 216 -22
rect 201 -25 205 -23
rect 207 -25 212 -23
rect 214 -25 216 -23
rect 201 -26 216 -25
rect 226 -23 234 -21
rect 226 -25 231 -23
rect 233 -25 234 -23
rect 210 -31 214 -26
rect 226 -27 234 -25
rect 257 -11 262 -6
rect 257 -13 258 -11
rect 260 -13 262 -11
rect 257 -15 262 -13
rect 210 -33 211 -31
rect 213 -33 214 -31
rect 210 -35 214 -33
rect 177 -39 183 -38
rect 177 -41 180 -39
rect 182 -41 183 -39
rect 177 -42 183 -41
rect 258 -31 262 -15
rect 267 -6 271 -5
rect 267 -8 268 -6
rect 270 -8 271 -6
rect 267 -14 271 -8
rect 267 -16 288 -14
rect 267 -18 272 -16
rect 274 -18 288 -16
rect 258 -33 259 -31
rect 261 -33 262 -31
rect 258 -37 262 -33
rect 267 -23 288 -22
rect 267 -25 268 -23
rect 270 -25 282 -23
rect 284 -25 288 -23
rect 267 -26 288 -25
rect 301 -4 303 -2
rect 299 -9 303 -4
rect 301 -11 303 -9
rect 267 -35 271 -26
rect 299 -27 303 -11
rect 315 -14 319 -5
rect 566 2 570 3
rect 557 -2 570 2
rect 355 -4 360 -2
rect 346 -6 351 -4
rect 315 -15 328 -14
rect 315 -17 320 -15
rect 322 -17 328 -15
rect 315 -18 328 -17
rect 299 -29 300 -27
rect 302 -29 303 -27
rect 299 -30 303 -29
rect 298 -32 303 -30
rect 298 -34 299 -32
rect 301 -34 303 -32
rect 298 -36 303 -34
rect 322 -23 336 -22
rect 322 -25 330 -23
rect 332 -25 336 -23
rect 322 -26 336 -25
rect 346 -8 347 -6
rect 349 -8 351 -6
rect 346 -13 351 -8
rect 346 -15 347 -13
rect 349 -15 351 -13
rect 346 -17 351 -15
rect 322 -29 327 -26
rect 322 -31 324 -29
rect 326 -31 327 -29
rect 322 -35 327 -31
rect 347 -23 351 -17
rect 347 -25 348 -23
rect 350 -25 351 -23
rect 257 -39 262 -37
rect 347 -37 351 -25
rect 257 -41 258 -39
rect 260 -41 262 -39
rect 257 -43 262 -41
rect 339 -39 347 -37
rect 349 -39 351 -37
rect 339 -43 351 -39
rect 355 -6 357 -4
rect 359 -6 360 -4
rect 355 -11 360 -6
rect 355 -13 357 -11
rect 359 -13 360 -11
rect 355 -15 360 -13
rect 355 -31 359 -15
rect 386 -15 424 -14
rect 386 -17 388 -15
rect 390 -17 424 -15
rect 386 -18 424 -17
rect 386 -21 391 -18
rect 383 -23 391 -21
rect 383 -25 384 -23
rect 386 -25 391 -23
rect 383 -27 391 -25
rect 401 -23 416 -22
rect 401 -25 403 -23
rect 405 -25 406 -23
rect 408 -25 410 -23
rect 412 -25 416 -23
rect 401 -26 416 -25
rect 355 -33 356 -31
rect 358 -33 359 -31
rect 355 -37 359 -33
rect 355 -39 360 -37
rect 403 -35 407 -26
rect 434 -7 440 -5
rect 434 -9 435 -7
rect 437 -9 440 -7
rect 434 -14 440 -9
rect 434 -16 435 -14
rect 437 -16 440 -14
rect 434 -18 440 -16
rect 436 -23 440 -18
rect 436 -25 437 -23
rect 439 -25 440 -23
rect 436 -38 440 -25
rect 355 -41 357 -39
rect 359 -41 360 -39
rect 355 -43 360 -41
rect 434 -39 440 -38
rect 434 -41 435 -39
rect 437 -41 440 -39
rect 434 -42 440 -41
rect 444 -7 450 -5
rect 524 -4 529 -2
rect 524 -6 525 -4
rect 527 -6 529 -4
rect 444 -9 447 -7
rect 449 -9 450 -7
rect 444 -10 450 -9
rect 444 -12 447 -10
rect 449 -12 450 -10
rect 444 -14 450 -12
rect 444 -16 447 -14
rect 449 -16 450 -14
rect 444 -18 450 -16
rect 444 -38 448 -18
rect 460 -15 498 -14
rect 460 -17 494 -15
rect 496 -17 498 -15
rect 460 -18 498 -17
rect 493 -21 498 -18
rect 468 -23 483 -22
rect 468 -25 472 -23
rect 474 -25 479 -23
rect 481 -25 483 -23
rect 468 -26 483 -25
rect 493 -23 501 -21
rect 493 -25 498 -23
rect 500 -25 501 -23
rect 477 -31 481 -26
rect 493 -27 501 -25
rect 524 -11 529 -6
rect 524 -13 525 -11
rect 527 -13 529 -11
rect 524 -15 529 -13
rect 477 -33 478 -31
rect 480 -33 481 -31
rect 477 -35 481 -33
rect 444 -39 450 -38
rect 444 -41 447 -39
rect 449 -41 450 -39
rect 444 -42 450 -41
rect 525 -31 529 -15
rect 534 -6 538 -5
rect 534 -8 535 -6
rect 537 -8 538 -6
rect 534 -14 538 -8
rect 534 -16 555 -14
rect 534 -18 539 -16
rect 541 -18 555 -16
rect 525 -33 526 -31
rect 528 -33 529 -31
rect 525 -37 529 -33
rect 534 -23 555 -22
rect 534 -25 535 -23
rect 537 -25 549 -23
rect 551 -25 555 -23
rect 534 -26 555 -25
rect 568 -4 570 -2
rect 566 -9 570 -4
rect 568 -11 570 -9
rect 534 -35 538 -26
rect 566 -27 570 -11
rect 582 -14 586 -5
rect 833 2 837 3
rect 824 -2 837 2
rect 622 -4 627 -2
rect 613 -6 618 -4
rect 582 -15 595 -14
rect 582 -17 587 -15
rect 589 -17 595 -15
rect 582 -18 595 -17
rect 566 -29 567 -27
rect 569 -29 570 -27
rect 566 -30 570 -29
rect 565 -32 570 -30
rect 565 -34 566 -32
rect 568 -34 570 -32
rect 565 -36 570 -34
rect 589 -23 603 -22
rect 589 -25 597 -23
rect 599 -25 603 -23
rect 589 -26 603 -25
rect 613 -8 614 -6
rect 616 -8 618 -6
rect 613 -13 618 -8
rect 613 -15 614 -13
rect 616 -15 618 -13
rect 613 -17 618 -15
rect 589 -29 594 -26
rect 589 -31 591 -29
rect 593 -31 594 -29
rect 589 -35 594 -31
rect 614 -23 618 -17
rect 614 -25 615 -23
rect 617 -25 618 -23
rect 524 -39 529 -37
rect 614 -37 618 -25
rect 524 -41 525 -39
rect 527 -41 529 -39
rect 524 -43 529 -41
rect 606 -39 614 -37
rect 616 -39 618 -37
rect 606 -43 618 -39
rect 622 -6 624 -4
rect 626 -6 627 -4
rect 622 -11 627 -6
rect 622 -13 624 -11
rect 626 -13 627 -11
rect 622 -15 627 -13
rect 622 -31 626 -15
rect 653 -15 691 -14
rect 653 -17 655 -15
rect 657 -17 691 -15
rect 653 -18 691 -17
rect 653 -21 658 -18
rect 650 -23 658 -21
rect 650 -25 651 -23
rect 653 -25 658 -23
rect 650 -27 658 -25
rect 668 -23 683 -22
rect 668 -25 670 -23
rect 672 -25 673 -23
rect 675 -25 677 -23
rect 679 -25 683 -23
rect 668 -26 683 -25
rect 622 -33 623 -31
rect 625 -33 626 -31
rect 622 -37 626 -33
rect 622 -39 627 -37
rect 670 -35 674 -26
rect 701 -7 707 -5
rect 701 -9 702 -7
rect 704 -9 707 -7
rect 701 -14 707 -9
rect 701 -16 702 -14
rect 704 -16 707 -14
rect 701 -18 707 -16
rect 703 -23 707 -18
rect 703 -25 704 -23
rect 706 -25 707 -23
rect 703 -38 707 -25
rect 622 -41 624 -39
rect 626 -41 627 -39
rect 622 -43 627 -41
rect 701 -39 707 -38
rect 701 -41 702 -39
rect 704 -41 707 -39
rect 701 -42 707 -41
rect 711 -7 717 -5
rect 791 -4 796 -2
rect 791 -6 792 -4
rect 794 -6 796 -4
rect 711 -9 714 -7
rect 716 -9 717 -7
rect 711 -10 717 -9
rect 711 -12 714 -10
rect 716 -12 717 -10
rect 711 -14 717 -12
rect 711 -16 714 -14
rect 716 -16 717 -14
rect 711 -18 717 -16
rect 711 -38 715 -18
rect 727 -15 765 -14
rect 727 -17 761 -15
rect 763 -17 765 -15
rect 727 -18 765 -17
rect 760 -21 765 -18
rect 735 -23 750 -22
rect 735 -25 739 -23
rect 741 -25 746 -23
rect 748 -25 750 -23
rect 735 -26 750 -25
rect 760 -23 768 -21
rect 760 -25 765 -23
rect 767 -25 768 -23
rect 744 -31 748 -26
rect 760 -27 768 -25
rect 791 -11 796 -6
rect 791 -13 792 -11
rect 794 -13 796 -11
rect 791 -15 796 -13
rect 744 -33 745 -31
rect 747 -33 748 -31
rect 744 -35 748 -33
rect 711 -39 717 -38
rect 711 -41 714 -39
rect 716 -41 717 -39
rect 711 -42 717 -41
rect 792 -31 796 -15
rect 801 -6 805 -5
rect 801 -8 802 -6
rect 804 -8 805 -6
rect 801 -14 805 -8
rect 801 -16 822 -14
rect 801 -18 806 -16
rect 808 -18 822 -16
rect 792 -33 793 -31
rect 795 -33 796 -31
rect 792 -37 796 -33
rect 801 -23 822 -22
rect 801 -25 802 -23
rect 804 -25 816 -23
rect 818 -25 822 -23
rect 801 -26 822 -25
rect 835 -4 837 -2
rect 833 -9 837 -4
rect 835 -11 837 -9
rect 801 -35 805 -26
rect 833 -27 837 -11
rect 849 -14 853 -5
rect 1100 2 1104 3
rect 1091 -2 1104 2
rect 889 -4 894 -2
rect 880 -6 885 -4
rect 849 -15 862 -14
rect 849 -17 854 -15
rect 856 -17 862 -15
rect 849 -18 862 -17
rect 833 -29 834 -27
rect 836 -29 837 -27
rect 833 -30 837 -29
rect 832 -32 837 -30
rect 832 -34 833 -32
rect 835 -34 837 -32
rect 832 -36 837 -34
rect 856 -23 870 -22
rect 856 -25 864 -23
rect 866 -25 870 -23
rect 856 -26 870 -25
rect 880 -8 881 -6
rect 883 -8 885 -6
rect 880 -13 885 -8
rect 880 -15 881 -13
rect 883 -15 885 -13
rect 880 -17 885 -15
rect 856 -29 861 -26
rect 856 -31 858 -29
rect 860 -31 861 -29
rect 856 -35 861 -31
rect 881 -23 885 -17
rect 881 -25 882 -23
rect 884 -25 885 -23
rect 791 -39 796 -37
rect 881 -37 885 -25
rect 791 -41 792 -39
rect 794 -41 796 -39
rect 791 -43 796 -41
rect 873 -39 881 -37
rect 883 -39 885 -37
rect 873 -43 885 -39
rect 889 -6 891 -4
rect 893 -6 894 -4
rect 889 -11 894 -6
rect 889 -13 891 -11
rect 893 -13 894 -11
rect 889 -15 894 -13
rect 889 -31 893 -15
rect 920 -15 958 -14
rect 920 -17 922 -15
rect 924 -17 958 -15
rect 920 -18 958 -17
rect 920 -21 925 -18
rect 917 -23 925 -21
rect 917 -25 918 -23
rect 920 -25 925 -23
rect 917 -27 925 -25
rect 935 -23 950 -22
rect 935 -25 937 -23
rect 939 -25 940 -23
rect 942 -25 944 -23
rect 946 -25 950 -23
rect 935 -26 950 -25
rect 889 -33 890 -31
rect 892 -33 893 -31
rect 889 -37 893 -33
rect 889 -39 894 -37
rect 937 -35 941 -26
rect 968 -7 974 -5
rect 968 -9 969 -7
rect 971 -9 974 -7
rect 968 -14 974 -9
rect 968 -16 969 -14
rect 971 -16 974 -14
rect 968 -18 974 -16
rect 970 -23 974 -18
rect 970 -25 971 -23
rect 973 -25 974 -23
rect 970 -38 974 -25
rect 889 -41 891 -39
rect 893 -41 894 -39
rect 889 -43 894 -41
rect 968 -39 974 -38
rect 968 -41 969 -39
rect 971 -41 974 -39
rect 968 -42 974 -41
rect 978 -7 984 -5
rect 1058 -4 1063 -2
rect 1058 -6 1059 -4
rect 1061 -6 1063 -4
rect 978 -9 981 -7
rect 983 -9 984 -7
rect 978 -10 984 -9
rect 978 -12 981 -10
rect 983 -12 984 -10
rect 978 -14 984 -12
rect 978 -16 981 -14
rect 983 -16 984 -14
rect 978 -18 984 -16
rect 978 -38 982 -18
rect 994 -15 1032 -14
rect 994 -17 1028 -15
rect 1030 -17 1032 -15
rect 994 -18 1032 -17
rect 1027 -21 1032 -18
rect 1002 -23 1017 -22
rect 1002 -25 1006 -23
rect 1008 -25 1013 -23
rect 1015 -25 1017 -23
rect 1002 -26 1017 -25
rect 1027 -23 1035 -21
rect 1027 -25 1032 -23
rect 1034 -25 1035 -23
rect 1011 -31 1015 -26
rect 1027 -27 1035 -25
rect 1058 -11 1063 -6
rect 1058 -13 1059 -11
rect 1061 -13 1063 -11
rect 1058 -15 1063 -13
rect 1011 -33 1012 -31
rect 1014 -33 1015 -31
rect 1011 -35 1015 -33
rect 978 -39 984 -38
rect 978 -41 981 -39
rect 983 -41 984 -39
rect 978 -42 984 -41
rect 1059 -31 1063 -15
rect 1068 -6 1072 -5
rect 1068 -8 1069 -6
rect 1071 -8 1072 -6
rect 1068 -14 1072 -8
rect 1068 -16 1089 -14
rect 1068 -18 1073 -16
rect 1075 -18 1089 -16
rect 1059 -33 1060 -31
rect 1062 -33 1063 -31
rect 1059 -37 1063 -33
rect 1068 -23 1089 -22
rect 1068 -25 1069 -23
rect 1071 -25 1083 -23
rect 1085 -25 1089 -23
rect 1068 -26 1089 -25
rect 1102 -4 1104 -2
rect 1100 -9 1104 -4
rect 1102 -11 1104 -9
rect 1068 -35 1072 -26
rect 1100 -27 1104 -11
rect 1116 -14 1120 -5
rect 1367 2 1371 3
rect 1358 -2 1371 2
rect 1156 -4 1161 -2
rect 1147 -6 1152 -4
rect 1116 -15 1129 -14
rect 1116 -17 1121 -15
rect 1123 -17 1129 -15
rect 1116 -18 1129 -17
rect 1100 -29 1101 -27
rect 1103 -29 1104 -27
rect 1100 -30 1104 -29
rect 1099 -32 1104 -30
rect 1099 -34 1100 -32
rect 1102 -34 1104 -32
rect 1099 -36 1104 -34
rect 1123 -23 1137 -22
rect 1123 -25 1131 -23
rect 1133 -25 1137 -23
rect 1123 -26 1137 -25
rect 1147 -8 1148 -6
rect 1150 -8 1152 -6
rect 1147 -13 1152 -8
rect 1147 -15 1148 -13
rect 1150 -15 1152 -13
rect 1147 -17 1152 -15
rect 1123 -29 1128 -26
rect 1123 -31 1125 -29
rect 1127 -31 1128 -29
rect 1123 -35 1128 -31
rect 1148 -23 1152 -17
rect 1148 -25 1149 -23
rect 1151 -25 1152 -23
rect 1058 -39 1063 -37
rect 1148 -37 1152 -25
rect 1058 -41 1059 -39
rect 1061 -41 1063 -39
rect 1058 -43 1063 -41
rect 1140 -39 1148 -37
rect 1150 -39 1152 -37
rect 1140 -43 1152 -39
rect 1156 -6 1158 -4
rect 1160 -6 1161 -4
rect 1156 -11 1161 -6
rect 1156 -13 1158 -11
rect 1160 -13 1161 -11
rect 1156 -15 1161 -13
rect 1156 -31 1160 -15
rect 1187 -15 1225 -14
rect 1187 -17 1189 -15
rect 1191 -17 1225 -15
rect 1187 -18 1225 -17
rect 1187 -21 1192 -18
rect 1184 -23 1192 -21
rect 1184 -25 1185 -23
rect 1187 -25 1192 -23
rect 1184 -27 1192 -25
rect 1202 -23 1217 -22
rect 1202 -25 1204 -23
rect 1206 -25 1207 -23
rect 1209 -25 1211 -23
rect 1213 -25 1217 -23
rect 1202 -26 1217 -25
rect 1156 -33 1157 -31
rect 1159 -33 1160 -31
rect 1156 -37 1160 -33
rect 1156 -39 1161 -37
rect 1204 -35 1208 -26
rect 1235 -7 1241 -5
rect 1235 -9 1236 -7
rect 1238 -9 1241 -7
rect 1235 -14 1241 -9
rect 1235 -16 1236 -14
rect 1238 -16 1241 -14
rect 1235 -18 1241 -16
rect 1237 -23 1241 -18
rect 1237 -25 1238 -23
rect 1240 -25 1241 -23
rect 1237 -38 1241 -25
rect 1156 -41 1158 -39
rect 1160 -41 1161 -39
rect 1156 -43 1161 -41
rect 1235 -39 1241 -38
rect 1235 -41 1236 -39
rect 1238 -41 1241 -39
rect 1235 -42 1241 -41
rect 1245 -7 1251 -5
rect 1325 -4 1330 -2
rect 1325 -6 1326 -4
rect 1328 -6 1330 -4
rect 1245 -9 1248 -7
rect 1250 -9 1251 -7
rect 1245 -10 1251 -9
rect 1245 -12 1248 -10
rect 1250 -12 1251 -10
rect 1245 -14 1251 -12
rect 1245 -16 1248 -14
rect 1250 -16 1251 -14
rect 1245 -18 1251 -16
rect 1245 -38 1249 -18
rect 1261 -15 1299 -14
rect 1261 -17 1295 -15
rect 1297 -17 1299 -15
rect 1261 -18 1299 -17
rect 1294 -21 1299 -18
rect 1269 -23 1284 -22
rect 1269 -25 1273 -23
rect 1275 -25 1280 -23
rect 1282 -25 1284 -23
rect 1269 -26 1284 -25
rect 1294 -23 1302 -21
rect 1294 -25 1299 -23
rect 1301 -25 1302 -23
rect 1278 -31 1282 -26
rect 1294 -27 1302 -25
rect 1325 -11 1330 -6
rect 1325 -13 1326 -11
rect 1328 -13 1330 -11
rect 1325 -15 1330 -13
rect 1278 -33 1279 -31
rect 1281 -33 1282 -31
rect 1278 -35 1282 -33
rect 1245 -39 1251 -38
rect 1245 -41 1248 -39
rect 1250 -41 1251 -39
rect 1245 -42 1251 -41
rect 1326 -31 1330 -15
rect 1335 -6 1339 -5
rect 1335 -8 1336 -6
rect 1338 -8 1339 -6
rect 1335 -14 1339 -8
rect 1335 -16 1356 -14
rect 1335 -18 1340 -16
rect 1342 -18 1356 -16
rect 1326 -33 1327 -31
rect 1329 -33 1330 -31
rect 1326 -37 1330 -33
rect 1335 -23 1356 -22
rect 1335 -25 1336 -23
rect 1338 -25 1350 -23
rect 1352 -25 1356 -23
rect 1335 -26 1356 -25
rect 1369 -4 1371 -2
rect 1367 -9 1371 -4
rect 1369 -11 1371 -9
rect 1335 -35 1339 -26
rect 1367 -27 1371 -11
rect 1383 -14 1387 -5
rect 1634 2 1638 3
rect 1625 -2 1638 2
rect 1423 -4 1428 -2
rect 1414 -6 1419 -4
rect 1383 -15 1396 -14
rect 1383 -17 1388 -15
rect 1390 -17 1396 -15
rect 1383 -18 1396 -17
rect 1367 -29 1368 -27
rect 1370 -29 1371 -27
rect 1367 -30 1371 -29
rect 1366 -32 1371 -30
rect 1366 -34 1367 -32
rect 1369 -34 1371 -32
rect 1366 -36 1371 -34
rect 1390 -23 1404 -22
rect 1390 -25 1398 -23
rect 1400 -25 1404 -23
rect 1390 -26 1404 -25
rect 1414 -8 1415 -6
rect 1417 -8 1419 -6
rect 1414 -13 1419 -8
rect 1414 -15 1415 -13
rect 1417 -15 1419 -13
rect 1414 -17 1419 -15
rect 1390 -29 1395 -26
rect 1390 -31 1392 -29
rect 1394 -31 1395 -29
rect 1390 -35 1395 -31
rect 1415 -23 1419 -17
rect 1415 -25 1416 -23
rect 1418 -25 1419 -23
rect 1325 -39 1330 -37
rect 1415 -37 1419 -25
rect 1325 -41 1326 -39
rect 1328 -41 1330 -39
rect 1325 -43 1330 -41
rect 1407 -39 1415 -37
rect 1417 -39 1419 -37
rect 1407 -43 1419 -39
rect 1423 -6 1425 -4
rect 1427 -6 1428 -4
rect 1423 -11 1428 -6
rect 1423 -13 1425 -11
rect 1427 -13 1428 -11
rect 1423 -15 1428 -13
rect 1423 -31 1427 -15
rect 1454 -15 1492 -14
rect 1454 -17 1456 -15
rect 1458 -17 1492 -15
rect 1454 -18 1492 -17
rect 1454 -21 1459 -18
rect 1451 -23 1459 -21
rect 1451 -25 1452 -23
rect 1454 -25 1459 -23
rect 1451 -27 1459 -25
rect 1469 -23 1484 -22
rect 1469 -25 1471 -23
rect 1473 -25 1474 -23
rect 1476 -25 1478 -23
rect 1480 -25 1484 -23
rect 1469 -26 1484 -25
rect 1423 -33 1424 -31
rect 1426 -33 1427 -31
rect 1423 -37 1427 -33
rect 1423 -39 1428 -37
rect 1471 -35 1475 -26
rect 1502 -7 1508 -5
rect 1502 -9 1503 -7
rect 1505 -9 1508 -7
rect 1502 -14 1508 -9
rect 1502 -16 1503 -14
rect 1505 -16 1508 -14
rect 1502 -18 1508 -16
rect 1504 -23 1508 -18
rect 1504 -25 1505 -23
rect 1507 -25 1508 -23
rect 1504 -38 1508 -25
rect 1423 -41 1425 -39
rect 1427 -41 1428 -39
rect 1423 -43 1428 -41
rect 1502 -39 1508 -38
rect 1502 -41 1503 -39
rect 1505 -41 1508 -39
rect 1502 -42 1508 -41
rect 1512 -7 1518 -5
rect 1592 -4 1597 -2
rect 1592 -6 1593 -4
rect 1595 -6 1597 -4
rect 1512 -9 1515 -7
rect 1517 -9 1518 -7
rect 1512 -10 1518 -9
rect 1512 -12 1515 -10
rect 1517 -12 1518 -10
rect 1512 -14 1518 -12
rect 1512 -16 1515 -14
rect 1517 -16 1518 -14
rect 1512 -18 1518 -16
rect 1512 -38 1516 -18
rect 1528 -15 1566 -14
rect 1528 -17 1562 -15
rect 1564 -17 1566 -15
rect 1528 -18 1566 -17
rect 1561 -21 1566 -18
rect 1536 -23 1551 -22
rect 1536 -25 1540 -23
rect 1542 -25 1547 -23
rect 1549 -25 1551 -23
rect 1536 -26 1551 -25
rect 1561 -23 1569 -21
rect 1561 -25 1566 -23
rect 1568 -25 1569 -23
rect 1545 -31 1549 -26
rect 1561 -27 1569 -25
rect 1592 -11 1597 -6
rect 1592 -13 1593 -11
rect 1595 -13 1597 -11
rect 1592 -15 1597 -13
rect 1545 -33 1546 -31
rect 1548 -33 1549 -31
rect 1545 -35 1549 -33
rect 1512 -39 1518 -38
rect 1512 -41 1515 -39
rect 1517 -41 1518 -39
rect 1512 -42 1518 -41
rect 1593 -31 1597 -15
rect 1602 -6 1606 -5
rect 1602 -8 1603 -6
rect 1605 -8 1606 -6
rect 1602 -14 1606 -8
rect 1602 -16 1623 -14
rect 1602 -18 1607 -16
rect 1609 -18 1623 -16
rect 1593 -33 1594 -31
rect 1596 -33 1597 -31
rect 1593 -37 1597 -33
rect 1602 -23 1623 -22
rect 1602 -25 1603 -23
rect 1605 -25 1617 -23
rect 1619 -25 1623 -23
rect 1602 -26 1623 -25
rect 1636 -4 1638 -2
rect 1634 -9 1638 -4
rect 1636 -11 1638 -9
rect 1602 -35 1606 -26
rect 1634 -27 1638 -11
rect 1650 -14 1654 -5
rect 1901 2 1905 3
rect 1892 -2 1905 2
rect 1690 -4 1695 -2
rect 1681 -6 1686 -4
rect 1650 -15 1663 -14
rect 1650 -17 1655 -15
rect 1657 -17 1663 -15
rect 1650 -18 1663 -17
rect 1634 -29 1635 -27
rect 1637 -29 1638 -27
rect 1634 -30 1638 -29
rect 1633 -32 1638 -30
rect 1633 -34 1634 -32
rect 1636 -34 1638 -32
rect 1633 -36 1638 -34
rect 1657 -23 1671 -22
rect 1657 -25 1665 -23
rect 1667 -25 1671 -23
rect 1657 -26 1671 -25
rect 1681 -8 1682 -6
rect 1684 -8 1686 -6
rect 1681 -13 1686 -8
rect 1681 -15 1682 -13
rect 1684 -15 1686 -13
rect 1681 -17 1686 -15
rect 1657 -29 1662 -26
rect 1657 -31 1659 -29
rect 1661 -31 1662 -29
rect 1657 -35 1662 -31
rect 1682 -23 1686 -17
rect 1682 -25 1683 -23
rect 1685 -25 1686 -23
rect 1592 -39 1597 -37
rect 1682 -37 1686 -25
rect 1592 -41 1593 -39
rect 1595 -41 1597 -39
rect 1592 -43 1597 -41
rect 1674 -39 1682 -37
rect 1684 -39 1686 -37
rect 1674 -43 1686 -39
rect 1690 -6 1692 -4
rect 1694 -6 1695 -4
rect 1690 -11 1695 -6
rect 1690 -13 1692 -11
rect 1694 -13 1695 -11
rect 1690 -15 1695 -13
rect 1690 -31 1694 -15
rect 1721 -15 1759 -14
rect 1721 -17 1723 -15
rect 1725 -17 1759 -15
rect 1721 -18 1759 -17
rect 1721 -21 1726 -18
rect 1718 -23 1726 -21
rect 1718 -25 1719 -23
rect 1721 -25 1726 -23
rect 1718 -27 1726 -25
rect 1736 -23 1751 -22
rect 1736 -25 1738 -23
rect 1740 -25 1741 -23
rect 1743 -25 1745 -23
rect 1747 -25 1751 -23
rect 1736 -26 1751 -25
rect 1690 -33 1691 -31
rect 1693 -33 1694 -31
rect 1690 -37 1694 -33
rect 1690 -39 1695 -37
rect 1738 -35 1742 -26
rect 1769 -7 1775 -5
rect 1769 -9 1770 -7
rect 1772 -9 1775 -7
rect 1769 -14 1775 -9
rect 1769 -16 1770 -14
rect 1772 -16 1775 -14
rect 1769 -18 1775 -16
rect 1771 -23 1775 -18
rect 1771 -25 1772 -23
rect 1774 -25 1775 -23
rect 1771 -38 1775 -25
rect 1690 -41 1692 -39
rect 1694 -41 1695 -39
rect 1690 -43 1695 -41
rect 1769 -39 1775 -38
rect 1769 -41 1770 -39
rect 1772 -41 1775 -39
rect 1769 -42 1775 -41
rect 1779 -7 1785 -5
rect 1859 -4 1864 -2
rect 1859 -6 1860 -4
rect 1862 -6 1864 -4
rect 1779 -9 1782 -7
rect 1784 -9 1785 -7
rect 1779 -10 1785 -9
rect 1779 -12 1782 -10
rect 1784 -12 1785 -10
rect 1779 -14 1785 -12
rect 1779 -16 1782 -14
rect 1784 -16 1785 -14
rect 1779 -18 1785 -16
rect 1779 -38 1783 -18
rect 1795 -15 1833 -14
rect 1795 -17 1829 -15
rect 1831 -17 1833 -15
rect 1795 -18 1833 -17
rect 1828 -21 1833 -18
rect 1803 -23 1818 -22
rect 1803 -25 1807 -23
rect 1809 -25 1814 -23
rect 1816 -25 1818 -23
rect 1803 -26 1818 -25
rect 1828 -23 1836 -21
rect 1828 -25 1833 -23
rect 1835 -25 1836 -23
rect 1812 -31 1816 -26
rect 1828 -27 1836 -25
rect 1859 -11 1864 -6
rect 1859 -13 1860 -11
rect 1862 -13 1864 -11
rect 1859 -15 1864 -13
rect 1812 -33 1813 -31
rect 1815 -33 1816 -31
rect 1812 -35 1816 -33
rect 1779 -39 1785 -38
rect 1779 -41 1782 -39
rect 1784 -41 1785 -39
rect 1779 -42 1785 -41
rect 1860 -32 1864 -15
rect 1869 -6 1873 -5
rect 1869 -8 1870 -6
rect 1872 -8 1873 -6
rect 1869 -14 1873 -8
rect 1869 -16 1890 -14
rect 1869 -18 1874 -16
rect 1876 -18 1890 -16
rect 1860 -34 1861 -32
rect 1863 -34 1864 -32
rect 1860 -37 1864 -34
rect 1869 -23 1890 -22
rect 1869 -25 1870 -23
rect 1872 -25 1884 -23
rect 1886 -25 1890 -23
rect 1869 -26 1890 -25
rect 1903 -4 1905 -2
rect 1901 -9 1905 -4
rect 1903 -11 1905 -9
rect 1869 -35 1873 -26
rect 1901 -27 1905 -11
rect 1912 -3 1924 3
rect 1912 -15 1917 -3
rect 2187 2 2191 3
rect 2178 -2 2191 2
rect 1976 -4 1981 -2
rect 1912 -17 1914 -15
rect 1916 -17 1917 -15
rect 1912 -19 1917 -17
rect 1901 -29 1902 -27
rect 1904 -29 1905 -27
rect 1901 -30 1905 -29
rect 1900 -32 1905 -30
rect 1900 -34 1901 -32
rect 1903 -34 1905 -32
rect 1900 -36 1905 -34
rect 1928 -28 1933 -21
rect 1956 -6 1972 -5
rect 1956 -8 1958 -6
rect 1960 -8 1972 -6
rect 1956 -10 1972 -8
rect 1968 -15 1972 -10
rect 1968 -17 1969 -15
rect 1971 -17 1972 -15
rect 1928 -29 1930 -28
rect 1920 -30 1930 -29
rect 1932 -30 1933 -28
rect 1920 -32 1933 -30
rect 1920 -34 1925 -32
rect 1927 -34 1933 -32
rect 1920 -35 1933 -34
rect 1859 -39 1864 -37
rect 1968 -38 1972 -17
rect 1859 -41 1860 -39
rect 1862 -41 1864 -39
rect 1859 -43 1864 -41
rect 1948 -39 1972 -38
rect 1948 -41 1950 -39
rect 1952 -41 1972 -39
rect 1948 -42 1972 -41
rect 1976 -6 1978 -4
rect 1980 -6 1981 -4
rect 1976 -11 1981 -6
rect 1976 -13 1978 -11
rect 1980 -13 1981 -11
rect 1976 -15 1981 -13
rect 1976 -31 1980 -15
rect 2007 -15 2045 -14
rect 2007 -17 2018 -15
rect 2020 -17 2045 -15
rect 2007 -18 2045 -17
rect 2007 -21 2012 -18
rect 2004 -23 2012 -21
rect 2004 -25 2005 -23
rect 2007 -25 2012 -23
rect 2004 -27 2012 -25
rect 2022 -23 2037 -22
rect 2022 -25 2024 -23
rect 2026 -25 2031 -23
rect 2033 -25 2037 -23
rect 2022 -26 2037 -25
rect 1976 -33 1977 -31
rect 1979 -33 1980 -31
rect 1976 -37 1980 -33
rect 1976 -39 1981 -37
rect 2024 -35 2028 -26
rect 2055 -7 2061 -5
rect 2055 -9 2056 -7
rect 2058 -9 2061 -7
rect 2055 -14 2061 -9
rect 2055 -16 2056 -14
rect 2058 -16 2061 -14
rect 2055 -18 2061 -16
rect 2057 -23 2061 -18
rect 2057 -25 2058 -23
rect 2060 -25 2061 -23
rect 2057 -38 2061 -25
rect 1976 -41 1978 -39
rect 1980 -41 1981 -39
rect 1976 -43 1981 -41
rect 2055 -39 2061 -38
rect 2055 -41 2056 -39
rect 2058 -41 2061 -39
rect 2055 -42 2061 -41
rect 2065 -7 2071 -5
rect 2145 -4 2150 -2
rect 2145 -6 2146 -4
rect 2148 -6 2150 -4
rect 2065 -9 2068 -7
rect 2070 -9 2071 -7
rect 2065 -10 2071 -9
rect 2065 -12 2068 -10
rect 2070 -12 2071 -10
rect 2065 -14 2071 -12
rect 2065 -16 2068 -14
rect 2070 -16 2071 -14
rect 2065 -18 2071 -16
rect 2065 -38 2069 -18
rect 2081 -15 2119 -14
rect 2081 -17 2116 -15
rect 2118 -17 2119 -15
rect 2081 -18 2119 -17
rect 2114 -21 2119 -18
rect 2089 -23 2104 -22
rect 2089 -25 2093 -23
rect 2095 -25 2100 -23
rect 2102 -25 2104 -23
rect 2089 -26 2104 -25
rect 2114 -23 2122 -21
rect 2114 -25 2119 -23
rect 2121 -25 2122 -23
rect 2098 -31 2102 -26
rect 2114 -27 2122 -25
rect 2145 -11 2150 -6
rect 2145 -13 2146 -11
rect 2148 -13 2150 -11
rect 2145 -15 2150 -13
rect 2098 -33 2099 -31
rect 2101 -33 2102 -31
rect 2098 -35 2102 -33
rect 2065 -39 2071 -38
rect 2065 -41 2068 -39
rect 2070 -41 2071 -39
rect 2065 -42 2071 -41
rect 2146 -31 2150 -15
rect 2155 -6 2159 -5
rect 2155 -8 2156 -6
rect 2158 -8 2159 -6
rect 2155 -14 2159 -8
rect 2155 -16 2176 -14
rect 2155 -18 2160 -16
rect 2162 -18 2176 -16
rect 2146 -33 2147 -31
rect 2149 -33 2150 -31
rect 2146 -37 2150 -33
rect 2155 -23 2176 -22
rect 2155 -25 2156 -23
rect 2158 -25 2170 -23
rect 2172 -25 2176 -23
rect 2155 -26 2176 -25
rect 2189 -4 2191 -2
rect 2187 -9 2191 -4
rect 2189 -11 2191 -9
rect 2199 -3 2204 3
rect 2246 1 2259 2
rect 2246 -1 2255 1
rect 2257 -1 2259 1
rect 2199 -5 2201 -3
rect 2203 -5 2204 -3
rect 2246 -2 2259 -1
rect 2199 -6 2204 -5
rect 2199 -10 2212 -6
rect 2155 -35 2159 -26
rect 2187 -27 2191 -11
rect 2187 -29 2188 -27
rect 2190 -29 2191 -27
rect 2187 -30 2191 -29
rect 2186 -32 2191 -30
rect 2186 -34 2187 -32
rect 2189 -34 2191 -32
rect 2186 -36 2191 -34
rect 2145 -39 2150 -37
rect 2145 -41 2146 -39
rect 2148 -41 2150 -39
rect 2213 -23 2219 -21
rect 2213 -25 2214 -23
rect 2216 -25 2219 -23
rect 2213 -30 2219 -25
rect 2206 -31 2219 -30
rect 2206 -33 2210 -31
rect 2212 -33 2219 -31
rect 2231 -14 2243 -13
rect 2231 -16 2236 -14
rect 2238 -16 2243 -14
rect 2231 -18 2243 -16
rect 2231 -19 2241 -18
rect 2239 -20 2241 -19
rect 2239 -27 2243 -20
rect 2206 -34 2219 -33
rect 2255 -35 2259 -2
rect 2267 -3 2272 3
rect 2314 1 2327 2
rect 2314 -1 2323 1
rect 2325 -1 2327 1
rect 2267 -5 2269 -3
rect 2271 -5 2272 -3
rect 2314 -2 2327 -1
rect 2267 -6 2272 -5
rect 2267 -10 2280 -6
rect 2254 -37 2259 -35
rect 2145 -43 2150 -41
rect 2254 -39 2255 -37
rect 2257 -39 2259 -37
rect 2254 -41 2259 -39
rect 2281 -23 2287 -21
rect 2281 -25 2282 -23
rect 2284 -25 2287 -23
rect 2281 -30 2287 -25
rect 2274 -31 2287 -30
rect 2274 -33 2276 -31
rect 2278 -33 2287 -31
rect 2299 -14 2311 -13
rect 2299 -16 2300 -14
rect 2302 -16 2311 -14
rect 2299 -18 2311 -16
rect 2299 -19 2309 -18
rect 2307 -20 2309 -19
rect 2307 -27 2311 -20
rect 2274 -34 2287 -33
rect 2323 -35 2327 -2
rect 2322 -37 2327 -35
rect 2255 -43 2259 -41
rect 2322 -39 2323 -37
rect 2325 -39 2327 -37
rect 2322 -41 2327 -39
rect 2323 -43 2327 -41
rect 4 -49 2331 -48
rect 4 -51 29 -49
rect 31 -51 39 -49
rect 41 -51 69 -49
rect 71 -51 79 -49
rect 81 -51 298 -49
rect 300 -51 336 -49
rect 338 -51 346 -49
rect 348 -51 565 -49
rect 567 -51 603 -49
rect 605 -51 613 -49
rect 615 -51 832 -49
rect 834 -51 870 -49
rect 872 -51 880 -49
rect 882 -51 1099 -49
rect 1101 -51 1137 -49
rect 1139 -51 1147 -49
rect 1149 -51 1366 -49
rect 1368 -51 1404 -49
rect 1406 -51 1414 -49
rect 1416 -51 1633 -49
rect 1635 -51 1671 -49
rect 1673 -51 1681 -49
rect 1683 -51 1900 -49
rect 1902 -51 1915 -49
rect 1917 -51 1968 -49
rect 1970 -51 2186 -49
rect 2188 -51 2331 -49
rect 4 -55 2331 -51
rect 4 -57 2276 -55
rect 2278 -57 2331 -55
rect 4 -59 2331 -57
rect 4 -61 2311 -59
rect 2313 -61 2331 -59
rect 4 -63 29 -61
rect 31 -63 39 -61
rect 41 -63 69 -61
rect 71 -63 79 -61
rect 81 -63 298 -61
rect 300 -63 336 -61
rect 338 -63 346 -61
rect 348 -63 565 -61
rect 567 -63 603 -61
rect 605 -63 613 -61
rect 615 -63 832 -61
rect 834 -63 870 -61
rect 872 -63 880 -61
rect 882 -63 1099 -61
rect 1101 -63 1137 -61
rect 1139 -63 1147 -61
rect 1149 -63 1366 -61
rect 1368 -63 1404 -61
rect 1406 -63 1414 -61
rect 1416 -63 1633 -61
rect 1635 -63 1671 -61
rect 1673 -63 1681 -61
rect 1683 -63 1900 -61
rect 1902 -63 1915 -61
rect 1917 -63 1968 -61
rect 1970 -63 2186 -61
rect 2188 -63 2331 -61
rect 4 -64 2331 -63
rect 15 -83 20 -77
rect 32 -73 44 -69
rect 32 -75 40 -73
rect 42 -75 44 -73
rect 15 -85 17 -83
rect 19 -85 20 -83
rect 15 -86 20 -85
rect 15 -87 29 -86
rect 15 -89 23 -87
rect 25 -89 29 -87
rect 15 -90 29 -89
rect 8 -95 21 -94
rect 8 -97 13 -95
rect 15 -97 21 -95
rect 8 -98 21 -97
rect 8 -107 12 -98
rect 40 -95 44 -75
rect 55 -86 60 -77
rect 72 -73 84 -69
rect 72 -75 80 -73
rect 82 -75 84 -73
rect 55 -87 69 -86
rect 55 -89 63 -87
rect 65 -89 69 -87
rect 55 -90 69 -89
rect 39 -97 41 -95
rect 43 -97 44 -95
rect 39 -98 44 -97
rect 39 -100 40 -98
rect 42 -100 44 -98
rect 39 -106 44 -100
rect 39 -108 40 -106
rect 42 -108 44 -106
rect 48 -95 61 -94
rect 48 -97 53 -95
rect 55 -97 61 -95
rect 48 -98 61 -97
rect 48 -103 52 -98
rect 80 -87 84 -75
rect 80 -89 81 -87
rect 83 -89 84 -87
rect 80 -95 84 -89
rect 48 -105 49 -103
rect 51 -105 52 -103
rect 48 -107 52 -105
rect 79 -97 84 -95
rect 79 -99 80 -97
rect 82 -99 84 -97
rect 79 -104 84 -99
rect 39 -110 44 -108
rect 79 -106 80 -104
rect 82 -106 84 -104
rect 79 -108 84 -106
rect 88 -71 93 -69
rect 88 -73 90 -71
rect 92 -73 93 -71
rect 88 -75 93 -73
rect 88 -79 92 -75
rect 88 -81 89 -79
rect 91 -81 92 -79
rect 88 -97 92 -81
rect 167 -71 173 -70
rect 167 -73 168 -71
rect 170 -73 173 -71
rect 167 -74 173 -73
rect 88 -99 93 -97
rect 88 -101 90 -99
rect 92 -101 93 -99
rect 88 -106 93 -101
rect 116 -87 124 -85
rect 136 -86 140 -77
rect 116 -89 117 -87
rect 119 -89 124 -87
rect 116 -91 124 -89
rect 134 -87 149 -86
rect 134 -89 136 -87
rect 138 -89 139 -87
rect 141 -89 143 -87
rect 145 -89 149 -87
rect 134 -90 149 -89
rect 119 -94 124 -91
rect 169 -87 173 -74
rect 169 -89 170 -87
rect 172 -89 173 -87
rect 119 -95 157 -94
rect 119 -97 134 -95
rect 136 -97 157 -95
rect 119 -98 157 -97
rect 169 -94 173 -89
rect 167 -96 173 -94
rect 167 -98 168 -96
rect 170 -98 173 -96
rect 167 -103 173 -98
rect 167 -105 168 -103
rect 170 -105 173 -103
rect 88 -108 90 -106
rect 92 -108 93 -106
rect 88 -110 93 -108
rect 167 -107 173 -105
rect 177 -71 183 -70
rect 177 -73 180 -71
rect 182 -73 183 -71
rect 177 -74 183 -73
rect 257 -70 264 -69
rect 257 -71 261 -70
rect 257 -73 258 -71
rect 260 -72 261 -71
rect 263 -72 264 -70
rect 260 -73 264 -72
rect 177 -94 181 -74
rect 210 -79 214 -77
rect 210 -81 211 -79
rect 213 -81 214 -79
rect 177 -96 183 -94
rect 177 -98 180 -96
rect 182 -98 183 -96
rect 177 -100 183 -98
rect 177 -102 180 -100
rect 182 -102 183 -100
rect 177 -103 183 -102
rect 177 -105 180 -103
rect 182 -105 183 -103
rect 177 -107 183 -105
rect 210 -86 214 -81
rect 257 -75 264 -73
rect 201 -87 216 -86
rect 201 -89 205 -87
rect 207 -89 212 -87
rect 214 -89 216 -87
rect 201 -90 216 -89
rect 226 -87 234 -85
rect 226 -89 231 -87
rect 233 -89 234 -87
rect 226 -91 234 -89
rect 226 -92 231 -91
rect 226 -94 228 -92
rect 230 -94 231 -92
rect 193 -98 231 -94
rect 258 -97 262 -75
rect 267 -81 271 -80
rect 267 -83 268 -81
rect 270 -83 271 -81
rect 267 -86 271 -83
rect 267 -87 288 -86
rect 267 -89 282 -87
rect 284 -89 288 -87
rect 267 -90 288 -89
rect 298 -78 303 -76
rect 298 -80 299 -78
rect 301 -80 303 -78
rect 298 -82 303 -80
rect 257 -99 262 -97
rect 257 -101 258 -99
rect 260 -101 262 -99
rect 257 -106 262 -101
rect 257 -108 258 -106
rect 260 -108 262 -106
rect 267 -96 272 -94
rect 274 -96 288 -94
rect 267 -98 288 -96
rect 267 -100 271 -98
rect 267 -102 268 -100
rect 270 -102 271 -100
rect 267 -107 271 -102
rect 257 -110 262 -108
rect 299 -101 303 -82
rect 322 -86 327 -77
rect 339 -73 351 -69
rect 339 -75 347 -73
rect 349 -75 351 -73
rect 322 -87 336 -86
rect 322 -89 330 -87
rect 332 -89 336 -87
rect 322 -90 336 -89
rect 301 -103 303 -101
rect 299 -108 303 -103
rect 315 -95 328 -94
rect 315 -97 320 -95
rect 322 -97 328 -95
rect 315 -98 328 -97
rect 315 -103 319 -98
rect 347 -87 351 -75
rect 347 -89 348 -87
rect 350 -89 351 -87
rect 347 -95 351 -89
rect 315 -105 316 -103
rect 318 -105 319 -103
rect 315 -107 319 -105
rect 346 -97 351 -95
rect 346 -99 347 -97
rect 349 -99 351 -97
rect 346 -104 351 -99
rect 301 -110 303 -108
rect 290 -111 303 -110
rect 290 -113 292 -111
rect 294 -113 303 -111
rect 290 -114 303 -113
rect 299 -115 303 -114
rect 346 -106 347 -104
rect 349 -106 351 -104
rect 346 -108 351 -106
rect 355 -71 360 -69
rect 355 -73 357 -71
rect 359 -73 360 -71
rect 355 -75 360 -73
rect 355 -79 359 -75
rect 355 -81 356 -79
rect 358 -81 359 -79
rect 355 -97 359 -81
rect 434 -71 440 -70
rect 434 -73 435 -71
rect 437 -73 440 -71
rect 434 -74 440 -73
rect 355 -99 360 -97
rect 355 -101 357 -99
rect 359 -101 360 -99
rect 355 -106 360 -101
rect 383 -87 391 -85
rect 403 -86 407 -77
rect 383 -89 384 -87
rect 386 -89 391 -87
rect 383 -91 391 -89
rect 401 -87 416 -86
rect 401 -89 403 -87
rect 405 -89 406 -87
rect 408 -89 410 -87
rect 412 -89 416 -87
rect 401 -90 416 -89
rect 386 -94 391 -91
rect 436 -87 440 -74
rect 436 -89 437 -87
rect 439 -89 440 -87
rect 386 -95 424 -94
rect 386 -97 401 -95
rect 403 -97 424 -95
rect 386 -98 424 -97
rect 436 -94 440 -89
rect 434 -96 440 -94
rect 434 -98 435 -96
rect 437 -98 440 -96
rect 434 -103 440 -98
rect 434 -105 435 -103
rect 437 -105 440 -103
rect 355 -108 357 -106
rect 359 -108 360 -106
rect 355 -110 360 -108
rect 434 -107 440 -105
rect 444 -71 450 -70
rect 444 -73 447 -71
rect 449 -73 450 -71
rect 444 -74 450 -73
rect 524 -70 531 -69
rect 524 -71 528 -70
rect 524 -73 525 -71
rect 527 -72 528 -71
rect 530 -72 531 -70
rect 527 -73 531 -72
rect 444 -94 448 -74
rect 477 -79 481 -77
rect 477 -81 478 -79
rect 480 -81 481 -79
rect 444 -96 450 -94
rect 444 -98 447 -96
rect 449 -98 450 -96
rect 444 -100 450 -98
rect 444 -102 447 -100
rect 449 -102 450 -100
rect 444 -103 450 -102
rect 444 -105 447 -103
rect 449 -105 450 -103
rect 444 -107 450 -105
rect 477 -86 481 -81
rect 524 -75 531 -73
rect 468 -87 483 -86
rect 468 -89 472 -87
rect 474 -89 479 -87
rect 481 -89 483 -87
rect 468 -90 483 -89
rect 493 -87 501 -85
rect 493 -89 498 -87
rect 500 -89 501 -87
rect 493 -91 501 -89
rect 493 -92 498 -91
rect 493 -94 495 -92
rect 497 -94 498 -92
rect 460 -98 498 -94
rect 525 -97 529 -75
rect 534 -81 538 -80
rect 534 -83 535 -81
rect 537 -83 538 -81
rect 534 -86 538 -83
rect 534 -87 555 -86
rect 534 -89 549 -87
rect 551 -89 555 -87
rect 534 -90 555 -89
rect 565 -78 570 -76
rect 565 -80 566 -78
rect 568 -80 570 -78
rect 565 -82 570 -80
rect 524 -99 529 -97
rect 524 -101 525 -99
rect 527 -101 529 -99
rect 524 -106 529 -101
rect 524 -108 525 -106
rect 527 -108 529 -106
rect 534 -96 539 -94
rect 541 -96 555 -94
rect 534 -98 555 -96
rect 534 -100 538 -98
rect 534 -102 535 -100
rect 537 -102 538 -100
rect 534 -107 538 -102
rect 524 -110 529 -108
rect 566 -101 570 -82
rect 589 -86 594 -77
rect 606 -73 618 -69
rect 606 -75 614 -73
rect 616 -75 618 -73
rect 589 -87 603 -86
rect 589 -89 597 -87
rect 599 -89 603 -87
rect 589 -90 603 -89
rect 568 -103 570 -101
rect 566 -108 570 -103
rect 582 -95 595 -94
rect 582 -97 587 -95
rect 589 -97 595 -95
rect 582 -98 595 -97
rect 582 -103 586 -98
rect 614 -87 618 -75
rect 614 -89 615 -87
rect 617 -89 618 -87
rect 614 -95 618 -89
rect 582 -105 583 -103
rect 585 -105 586 -103
rect 582 -107 586 -105
rect 613 -97 618 -95
rect 613 -99 614 -97
rect 616 -99 618 -97
rect 613 -104 618 -99
rect 568 -110 570 -108
rect 557 -111 570 -110
rect 557 -113 559 -111
rect 561 -113 570 -111
rect 557 -114 570 -113
rect 566 -115 570 -114
rect 613 -106 614 -104
rect 616 -106 618 -104
rect 613 -108 618 -106
rect 622 -71 627 -69
rect 622 -73 624 -71
rect 626 -73 627 -71
rect 622 -75 627 -73
rect 622 -79 626 -75
rect 622 -81 623 -79
rect 625 -81 626 -79
rect 622 -97 626 -81
rect 701 -71 707 -70
rect 701 -73 702 -71
rect 704 -73 707 -71
rect 701 -74 707 -73
rect 622 -99 627 -97
rect 622 -101 624 -99
rect 626 -101 627 -99
rect 622 -106 627 -101
rect 650 -87 658 -85
rect 670 -86 674 -77
rect 650 -89 651 -87
rect 653 -89 658 -87
rect 650 -91 658 -89
rect 668 -87 683 -86
rect 668 -89 670 -87
rect 672 -89 673 -87
rect 675 -89 677 -87
rect 679 -89 683 -87
rect 668 -90 683 -89
rect 653 -94 658 -91
rect 703 -87 707 -74
rect 703 -89 704 -87
rect 706 -89 707 -87
rect 653 -95 691 -94
rect 653 -97 668 -95
rect 670 -97 691 -95
rect 653 -98 691 -97
rect 703 -94 707 -89
rect 701 -96 707 -94
rect 701 -98 702 -96
rect 704 -98 707 -96
rect 701 -103 707 -98
rect 701 -105 702 -103
rect 704 -105 707 -103
rect 622 -108 624 -106
rect 626 -108 627 -106
rect 622 -110 627 -108
rect 701 -107 707 -105
rect 711 -71 717 -70
rect 711 -73 714 -71
rect 716 -73 717 -71
rect 711 -74 717 -73
rect 791 -70 798 -69
rect 791 -71 795 -70
rect 791 -73 792 -71
rect 794 -72 795 -71
rect 797 -72 798 -70
rect 794 -73 798 -72
rect 711 -94 715 -74
rect 744 -79 748 -77
rect 744 -81 745 -79
rect 747 -81 748 -79
rect 711 -96 717 -94
rect 711 -98 714 -96
rect 716 -98 717 -96
rect 711 -100 717 -98
rect 711 -102 714 -100
rect 716 -102 717 -100
rect 711 -103 717 -102
rect 711 -105 714 -103
rect 716 -105 717 -103
rect 711 -107 717 -105
rect 744 -86 748 -81
rect 791 -75 798 -73
rect 735 -87 750 -86
rect 735 -89 739 -87
rect 741 -89 746 -87
rect 748 -89 750 -87
rect 735 -90 750 -89
rect 760 -87 768 -85
rect 760 -89 765 -87
rect 767 -89 768 -87
rect 760 -91 768 -89
rect 760 -92 765 -91
rect 760 -94 762 -92
rect 764 -94 765 -92
rect 727 -98 765 -94
rect 792 -97 796 -75
rect 801 -81 805 -80
rect 801 -83 802 -81
rect 804 -83 805 -81
rect 801 -86 805 -83
rect 801 -87 822 -86
rect 801 -89 816 -87
rect 818 -89 822 -87
rect 801 -90 822 -89
rect 832 -78 837 -76
rect 832 -80 833 -78
rect 835 -80 837 -78
rect 832 -82 837 -80
rect 791 -99 796 -97
rect 791 -101 792 -99
rect 794 -101 796 -99
rect 791 -106 796 -101
rect 791 -108 792 -106
rect 794 -108 796 -106
rect 801 -96 806 -94
rect 808 -96 822 -94
rect 801 -98 822 -96
rect 801 -100 805 -98
rect 801 -102 802 -100
rect 804 -102 805 -100
rect 801 -107 805 -102
rect 791 -110 796 -108
rect 833 -101 837 -82
rect 856 -86 861 -77
rect 873 -73 885 -69
rect 873 -75 881 -73
rect 883 -75 885 -73
rect 856 -87 870 -86
rect 856 -89 864 -87
rect 866 -89 870 -87
rect 856 -90 870 -89
rect 835 -103 837 -101
rect 833 -108 837 -103
rect 849 -95 862 -94
rect 849 -97 854 -95
rect 856 -97 862 -95
rect 849 -98 862 -97
rect 849 -103 853 -98
rect 881 -87 885 -75
rect 881 -89 882 -87
rect 884 -89 885 -87
rect 881 -95 885 -89
rect 849 -105 850 -103
rect 852 -105 853 -103
rect 849 -107 853 -105
rect 880 -97 885 -95
rect 880 -99 881 -97
rect 883 -99 885 -97
rect 880 -104 885 -99
rect 835 -110 837 -108
rect 824 -111 837 -110
rect 824 -113 826 -111
rect 828 -113 837 -111
rect 824 -114 837 -113
rect 833 -115 837 -114
rect 880 -106 881 -104
rect 883 -106 885 -104
rect 880 -108 885 -106
rect 889 -71 894 -69
rect 889 -73 891 -71
rect 893 -73 894 -71
rect 889 -75 894 -73
rect 889 -79 893 -75
rect 889 -81 890 -79
rect 892 -81 893 -79
rect 889 -97 893 -81
rect 968 -71 974 -70
rect 968 -73 969 -71
rect 971 -73 974 -71
rect 968 -74 974 -73
rect 889 -99 894 -97
rect 889 -101 891 -99
rect 893 -101 894 -99
rect 889 -106 894 -101
rect 917 -87 925 -85
rect 937 -86 941 -77
rect 917 -89 918 -87
rect 920 -89 925 -87
rect 917 -91 925 -89
rect 935 -87 950 -86
rect 935 -89 937 -87
rect 939 -89 940 -87
rect 942 -89 944 -87
rect 946 -89 950 -87
rect 935 -90 950 -89
rect 920 -94 925 -91
rect 970 -87 974 -74
rect 970 -89 971 -87
rect 973 -89 974 -87
rect 920 -95 958 -94
rect 920 -97 935 -95
rect 937 -97 958 -95
rect 920 -98 958 -97
rect 970 -94 974 -89
rect 968 -96 974 -94
rect 968 -98 969 -96
rect 971 -98 974 -96
rect 968 -103 974 -98
rect 968 -105 969 -103
rect 971 -105 974 -103
rect 889 -108 891 -106
rect 893 -108 894 -106
rect 889 -110 894 -108
rect 968 -107 974 -105
rect 978 -71 984 -70
rect 978 -73 981 -71
rect 983 -73 984 -71
rect 978 -74 984 -73
rect 1058 -70 1065 -69
rect 1058 -71 1062 -70
rect 1058 -73 1059 -71
rect 1061 -72 1062 -71
rect 1064 -72 1065 -70
rect 1061 -73 1065 -72
rect 978 -94 982 -74
rect 1011 -79 1015 -77
rect 1011 -81 1012 -79
rect 1014 -81 1015 -79
rect 978 -96 984 -94
rect 978 -98 981 -96
rect 983 -98 984 -96
rect 978 -100 984 -98
rect 978 -102 981 -100
rect 983 -102 984 -100
rect 978 -103 984 -102
rect 978 -105 981 -103
rect 983 -105 984 -103
rect 978 -107 984 -105
rect 1011 -86 1015 -81
rect 1058 -75 1065 -73
rect 1002 -87 1017 -86
rect 1002 -89 1006 -87
rect 1008 -89 1013 -87
rect 1015 -89 1017 -87
rect 1002 -90 1017 -89
rect 1027 -87 1035 -85
rect 1027 -89 1032 -87
rect 1034 -89 1035 -87
rect 1027 -91 1035 -89
rect 1027 -92 1032 -91
rect 1027 -94 1029 -92
rect 1031 -94 1032 -92
rect 994 -98 1032 -94
rect 1059 -97 1063 -75
rect 1068 -81 1072 -80
rect 1068 -83 1069 -81
rect 1071 -83 1072 -81
rect 1068 -86 1072 -83
rect 1068 -87 1089 -86
rect 1068 -89 1083 -87
rect 1085 -89 1089 -87
rect 1068 -90 1089 -89
rect 1099 -78 1104 -76
rect 1099 -80 1100 -78
rect 1102 -80 1104 -78
rect 1099 -82 1104 -80
rect 1058 -99 1063 -97
rect 1058 -101 1059 -99
rect 1061 -101 1063 -99
rect 1058 -106 1063 -101
rect 1058 -108 1059 -106
rect 1061 -108 1063 -106
rect 1068 -96 1073 -94
rect 1075 -96 1089 -94
rect 1068 -98 1089 -96
rect 1068 -100 1072 -98
rect 1068 -102 1069 -100
rect 1071 -102 1072 -100
rect 1068 -107 1072 -102
rect 1058 -110 1063 -108
rect 1100 -101 1104 -82
rect 1123 -86 1128 -77
rect 1140 -73 1152 -69
rect 1140 -75 1148 -73
rect 1150 -75 1152 -73
rect 1123 -87 1137 -86
rect 1123 -89 1131 -87
rect 1133 -89 1137 -87
rect 1123 -90 1137 -89
rect 1102 -103 1104 -101
rect 1100 -108 1104 -103
rect 1116 -95 1129 -94
rect 1116 -97 1121 -95
rect 1123 -97 1129 -95
rect 1116 -98 1129 -97
rect 1116 -103 1120 -98
rect 1148 -87 1152 -75
rect 1148 -89 1149 -87
rect 1151 -89 1152 -87
rect 1148 -95 1152 -89
rect 1116 -105 1117 -103
rect 1119 -105 1120 -103
rect 1116 -107 1120 -105
rect 1147 -97 1152 -95
rect 1147 -99 1148 -97
rect 1150 -99 1152 -97
rect 1147 -104 1152 -99
rect 1102 -110 1104 -108
rect 1091 -111 1104 -110
rect 1091 -113 1093 -111
rect 1095 -113 1104 -111
rect 1091 -114 1104 -113
rect 1100 -115 1104 -114
rect 1147 -106 1148 -104
rect 1150 -106 1152 -104
rect 1147 -108 1152 -106
rect 1156 -71 1161 -69
rect 1156 -73 1158 -71
rect 1160 -73 1161 -71
rect 1156 -75 1161 -73
rect 1156 -79 1160 -75
rect 1156 -81 1157 -79
rect 1159 -81 1160 -79
rect 1156 -97 1160 -81
rect 1235 -71 1241 -70
rect 1235 -73 1236 -71
rect 1238 -73 1241 -71
rect 1235 -74 1241 -73
rect 1156 -99 1161 -97
rect 1156 -101 1158 -99
rect 1160 -101 1161 -99
rect 1156 -106 1161 -101
rect 1184 -87 1192 -85
rect 1204 -86 1208 -77
rect 1184 -89 1185 -87
rect 1187 -89 1192 -87
rect 1184 -91 1192 -89
rect 1202 -87 1217 -86
rect 1202 -89 1204 -87
rect 1206 -89 1207 -87
rect 1209 -89 1211 -87
rect 1213 -89 1217 -87
rect 1202 -90 1217 -89
rect 1187 -94 1192 -91
rect 1237 -87 1241 -74
rect 1237 -89 1238 -87
rect 1240 -89 1241 -87
rect 1187 -95 1225 -94
rect 1187 -97 1202 -95
rect 1204 -97 1225 -95
rect 1187 -98 1225 -97
rect 1237 -94 1241 -89
rect 1235 -96 1241 -94
rect 1235 -98 1236 -96
rect 1238 -98 1241 -96
rect 1235 -103 1241 -98
rect 1235 -105 1236 -103
rect 1238 -105 1241 -103
rect 1156 -108 1158 -106
rect 1160 -108 1161 -106
rect 1156 -110 1161 -108
rect 1235 -107 1241 -105
rect 1245 -71 1251 -70
rect 1245 -73 1248 -71
rect 1250 -73 1251 -71
rect 1245 -74 1251 -73
rect 1325 -70 1332 -69
rect 1325 -71 1329 -70
rect 1325 -73 1326 -71
rect 1328 -72 1329 -71
rect 1331 -72 1332 -70
rect 1328 -73 1332 -72
rect 1245 -94 1249 -74
rect 1278 -79 1282 -77
rect 1278 -81 1279 -79
rect 1281 -81 1282 -79
rect 1245 -96 1251 -94
rect 1245 -98 1248 -96
rect 1250 -98 1251 -96
rect 1245 -100 1251 -98
rect 1245 -102 1248 -100
rect 1250 -102 1251 -100
rect 1245 -103 1251 -102
rect 1245 -105 1248 -103
rect 1250 -105 1251 -103
rect 1245 -107 1251 -105
rect 1278 -86 1282 -81
rect 1325 -75 1332 -73
rect 1269 -87 1284 -86
rect 1269 -89 1273 -87
rect 1275 -89 1280 -87
rect 1282 -89 1284 -87
rect 1269 -90 1284 -89
rect 1294 -87 1302 -85
rect 1294 -89 1299 -87
rect 1301 -89 1302 -87
rect 1294 -91 1302 -89
rect 1294 -92 1299 -91
rect 1294 -94 1296 -92
rect 1298 -94 1299 -92
rect 1261 -98 1299 -94
rect 1326 -97 1330 -75
rect 1335 -81 1339 -80
rect 1335 -83 1336 -81
rect 1338 -83 1339 -81
rect 1335 -86 1339 -83
rect 1335 -87 1356 -86
rect 1335 -89 1350 -87
rect 1352 -89 1356 -87
rect 1335 -90 1356 -89
rect 1366 -78 1371 -76
rect 1366 -80 1367 -78
rect 1369 -80 1371 -78
rect 1366 -82 1371 -80
rect 1325 -99 1330 -97
rect 1325 -101 1326 -99
rect 1328 -101 1330 -99
rect 1325 -106 1330 -101
rect 1325 -108 1326 -106
rect 1328 -108 1330 -106
rect 1335 -96 1340 -94
rect 1342 -96 1356 -94
rect 1335 -98 1356 -96
rect 1335 -100 1339 -98
rect 1335 -102 1336 -100
rect 1338 -102 1339 -100
rect 1335 -107 1339 -102
rect 1325 -110 1330 -108
rect 1367 -101 1371 -82
rect 1390 -86 1395 -77
rect 1407 -73 1419 -69
rect 1407 -75 1415 -73
rect 1417 -75 1419 -73
rect 1390 -87 1404 -86
rect 1390 -89 1398 -87
rect 1400 -89 1404 -87
rect 1390 -90 1404 -89
rect 1369 -103 1371 -101
rect 1367 -108 1371 -103
rect 1383 -95 1396 -94
rect 1383 -97 1388 -95
rect 1390 -97 1396 -95
rect 1383 -98 1396 -97
rect 1383 -103 1387 -98
rect 1415 -87 1419 -75
rect 1415 -89 1416 -87
rect 1418 -89 1419 -87
rect 1415 -95 1419 -89
rect 1383 -105 1384 -103
rect 1386 -105 1387 -103
rect 1383 -107 1387 -105
rect 1414 -97 1419 -95
rect 1414 -99 1415 -97
rect 1417 -99 1419 -97
rect 1414 -104 1419 -99
rect 1369 -110 1371 -108
rect 1358 -111 1371 -110
rect 1358 -113 1360 -111
rect 1362 -113 1371 -111
rect 1358 -114 1371 -113
rect 1367 -115 1371 -114
rect 1414 -106 1415 -104
rect 1417 -106 1419 -104
rect 1414 -108 1419 -106
rect 1423 -71 1428 -69
rect 1423 -73 1425 -71
rect 1427 -73 1428 -71
rect 1423 -75 1428 -73
rect 1423 -79 1427 -75
rect 1423 -81 1424 -79
rect 1426 -81 1427 -79
rect 1423 -97 1427 -81
rect 1502 -71 1508 -70
rect 1502 -73 1503 -71
rect 1505 -73 1508 -71
rect 1502 -74 1508 -73
rect 1423 -99 1428 -97
rect 1423 -101 1425 -99
rect 1427 -101 1428 -99
rect 1423 -106 1428 -101
rect 1451 -87 1459 -85
rect 1471 -86 1475 -77
rect 1451 -89 1452 -87
rect 1454 -89 1459 -87
rect 1451 -91 1459 -89
rect 1469 -87 1484 -86
rect 1469 -89 1471 -87
rect 1473 -89 1474 -87
rect 1476 -89 1478 -87
rect 1480 -89 1484 -87
rect 1469 -90 1484 -89
rect 1454 -94 1459 -91
rect 1504 -87 1508 -74
rect 1504 -89 1505 -87
rect 1507 -89 1508 -87
rect 1454 -95 1492 -94
rect 1454 -97 1469 -95
rect 1471 -97 1492 -95
rect 1454 -98 1492 -97
rect 1504 -94 1508 -89
rect 1502 -96 1508 -94
rect 1502 -98 1503 -96
rect 1505 -98 1508 -96
rect 1502 -103 1508 -98
rect 1502 -105 1503 -103
rect 1505 -105 1508 -103
rect 1423 -108 1425 -106
rect 1427 -108 1428 -106
rect 1423 -110 1428 -108
rect 1502 -107 1508 -105
rect 1512 -71 1518 -70
rect 1512 -73 1515 -71
rect 1517 -73 1518 -71
rect 1512 -74 1518 -73
rect 1592 -70 1599 -69
rect 1592 -71 1596 -70
rect 1592 -73 1593 -71
rect 1595 -72 1596 -71
rect 1598 -72 1599 -70
rect 1595 -73 1599 -72
rect 1512 -94 1516 -74
rect 1545 -79 1549 -77
rect 1545 -81 1546 -79
rect 1548 -81 1549 -79
rect 1512 -96 1518 -94
rect 1512 -98 1515 -96
rect 1517 -98 1518 -96
rect 1512 -100 1518 -98
rect 1512 -102 1515 -100
rect 1517 -102 1518 -100
rect 1512 -103 1518 -102
rect 1512 -105 1515 -103
rect 1517 -105 1518 -103
rect 1512 -107 1518 -105
rect 1545 -86 1549 -81
rect 1592 -75 1599 -73
rect 1536 -87 1551 -86
rect 1536 -89 1540 -87
rect 1542 -89 1547 -87
rect 1549 -89 1551 -87
rect 1536 -90 1551 -89
rect 1561 -87 1569 -85
rect 1561 -89 1566 -87
rect 1568 -89 1569 -87
rect 1561 -91 1569 -89
rect 1561 -92 1566 -91
rect 1561 -94 1563 -92
rect 1565 -94 1566 -92
rect 1528 -98 1566 -94
rect 1593 -97 1597 -75
rect 1602 -81 1606 -80
rect 1602 -83 1603 -81
rect 1605 -83 1606 -81
rect 1602 -86 1606 -83
rect 1602 -87 1623 -86
rect 1602 -89 1617 -87
rect 1619 -89 1623 -87
rect 1602 -90 1623 -89
rect 1633 -78 1638 -76
rect 1633 -80 1634 -78
rect 1636 -80 1638 -78
rect 1633 -82 1638 -80
rect 1592 -99 1597 -97
rect 1592 -101 1593 -99
rect 1595 -101 1597 -99
rect 1592 -106 1597 -101
rect 1592 -108 1593 -106
rect 1595 -108 1597 -106
rect 1602 -96 1607 -94
rect 1609 -96 1623 -94
rect 1602 -98 1623 -96
rect 1602 -100 1606 -98
rect 1602 -102 1603 -100
rect 1605 -102 1606 -100
rect 1602 -107 1606 -102
rect 1592 -110 1597 -108
rect 1634 -101 1638 -82
rect 1657 -86 1662 -77
rect 1674 -73 1686 -69
rect 1674 -75 1682 -73
rect 1684 -75 1686 -73
rect 1657 -87 1671 -86
rect 1657 -89 1665 -87
rect 1667 -89 1671 -87
rect 1657 -90 1671 -89
rect 1636 -103 1638 -101
rect 1634 -108 1638 -103
rect 1650 -95 1663 -94
rect 1650 -97 1655 -95
rect 1657 -97 1663 -95
rect 1650 -98 1663 -97
rect 1650 -103 1654 -98
rect 1682 -87 1686 -75
rect 1682 -89 1683 -87
rect 1685 -89 1686 -87
rect 1682 -95 1686 -89
rect 1650 -105 1651 -103
rect 1653 -105 1654 -103
rect 1650 -107 1654 -105
rect 1681 -97 1686 -95
rect 1681 -99 1682 -97
rect 1684 -99 1686 -97
rect 1681 -104 1686 -99
rect 1636 -110 1638 -108
rect 1625 -111 1638 -110
rect 1625 -113 1627 -111
rect 1629 -113 1638 -111
rect 1625 -114 1638 -113
rect 1634 -115 1638 -114
rect 1681 -106 1682 -104
rect 1684 -106 1686 -104
rect 1681 -108 1686 -106
rect 1690 -71 1695 -69
rect 1690 -73 1692 -71
rect 1694 -73 1695 -71
rect 1690 -75 1695 -73
rect 1690 -79 1694 -75
rect 1690 -81 1691 -79
rect 1693 -81 1694 -79
rect 1690 -97 1694 -81
rect 1769 -71 1775 -70
rect 1769 -73 1770 -71
rect 1772 -73 1775 -71
rect 1769 -74 1775 -73
rect 1690 -99 1695 -97
rect 1690 -101 1692 -99
rect 1694 -101 1695 -99
rect 1690 -106 1695 -101
rect 1718 -87 1726 -85
rect 1738 -86 1742 -77
rect 1718 -89 1719 -87
rect 1721 -89 1726 -87
rect 1718 -91 1726 -89
rect 1736 -87 1751 -86
rect 1736 -89 1738 -87
rect 1740 -89 1741 -87
rect 1743 -89 1745 -87
rect 1747 -89 1751 -87
rect 1736 -90 1751 -89
rect 1721 -94 1726 -91
rect 1771 -87 1775 -74
rect 1771 -89 1772 -87
rect 1774 -89 1775 -87
rect 1721 -95 1759 -94
rect 1721 -97 1736 -95
rect 1738 -97 1759 -95
rect 1721 -98 1759 -97
rect 1771 -94 1775 -89
rect 1769 -96 1775 -94
rect 1769 -98 1770 -96
rect 1772 -98 1775 -96
rect 1769 -103 1775 -98
rect 1769 -105 1770 -103
rect 1772 -105 1775 -103
rect 1690 -108 1692 -106
rect 1694 -108 1695 -106
rect 1690 -110 1695 -108
rect 1769 -107 1775 -105
rect 1779 -71 1785 -70
rect 1779 -73 1782 -71
rect 1784 -73 1785 -71
rect 1779 -74 1785 -73
rect 1859 -70 1866 -69
rect 1859 -71 1863 -70
rect 1859 -73 1860 -71
rect 1862 -72 1863 -71
rect 1865 -72 1866 -70
rect 1862 -73 1866 -72
rect 1948 -71 1972 -70
rect 1779 -94 1783 -74
rect 1812 -79 1816 -77
rect 1812 -81 1813 -79
rect 1815 -81 1816 -79
rect 1779 -96 1785 -94
rect 1779 -98 1782 -96
rect 1784 -98 1785 -96
rect 1779 -100 1785 -98
rect 1779 -102 1782 -100
rect 1784 -102 1785 -100
rect 1779 -103 1785 -102
rect 1779 -105 1782 -103
rect 1784 -105 1785 -103
rect 1779 -107 1785 -105
rect 1812 -86 1816 -81
rect 1859 -75 1866 -73
rect 1948 -73 1950 -71
rect 1952 -73 1972 -71
rect 1948 -74 1972 -73
rect 1803 -87 1818 -86
rect 1803 -89 1807 -87
rect 1809 -89 1814 -87
rect 1816 -89 1818 -87
rect 1803 -90 1818 -89
rect 1828 -87 1836 -85
rect 1828 -89 1833 -87
rect 1835 -89 1836 -87
rect 1828 -91 1836 -89
rect 1828 -92 1833 -91
rect 1828 -94 1830 -92
rect 1832 -94 1833 -92
rect 1795 -98 1833 -94
rect 1860 -97 1864 -75
rect 1869 -81 1873 -80
rect 1869 -83 1870 -81
rect 1872 -83 1873 -81
rect 1869 -86 1873 -83
rect 1869 -87 1890 -86
rect 1869 -89 1884 -87
rect 1886 -89 1890 -87
rect 1869 -90 1890 -89
rect 1900 -78 1905 -76
rect 1900 -80 1901 -78
rect 1903 -80 1905 -78
rect 1900 -82 1905 -80
rect 1859 -99 1864 -97
rect 1859 -101 1860 -99
rect 1862 -101 1864 -99
rect 1859 -106 1864 -101
rect 1859 -108 1860 -106
rect 1862 -108 1864 -106
rect 1869 -96 1874 -94
rect 1876 -96 1890 -94
rect 1869 -98 1890 -96
rect 1869 -100 1873 -98
rect 1869 -102 1870 -100
rect 1872 -102 1873 -100
rect 1869 -107 1873 -102
rect 1859 -110 1864 -108
rect 1901 -101 1905 -82
rect 1920 -78 1933 -77
rect 1920 -80 1925 -78
rect 1927 -80 1933 -78
rect 1920 -82 1933 -80
rect 1920 -83 1930 -82
rect 1928 -84 1930 -83
rect 1932 -84 1933 -82
rect 1903 -103 1905 -101
rect 1901 -108 1905 -103
rect 1903 -110 1905 -108
rect 1892 -111 1905 -110
rect 1892 -113 1894 -111
rect 1896 -113 1905 -111
rect 1892 -114 1905 -113
rect 1901 -115 1905 -114
rect 1912 -95 1917 -93
rect 1912 -97 1914 -95
rect 1916 -97 1917 -95
rect 1912 -109 1917 -97
rect 1928 -91 1933 -84
rect 1912 -115 1924 -109
rect 1968 -95 1972 -74
rect 1968 -97 1969 -95
rect 1971 -97 1972 -95
rect 1968 -102 1972 -97
rect 1956 -104 1972 -102
rect 1956 -106 1958 -104
rect 1960 -106 1972 -104
rect 1956 -107 1972 -106
rect 1976 -71 1981 -69
rect 1976 -73 1978 -71
rect 1980 -73 1981 -71
rect 1976 -75 1981 -73
rect 1976 -79 1980 -75
rect 1976 -81 1977 -79
rect 1979 -81 1980 -79
rect 1976 -97 1980 -81
rect 2055 -71 2061 -70
rect 2055 -73 2056 -71
rect 2058 -73 2061 -71
rect 2055 -74 2061 -73
rect 1976 -99 1981 -97
rect 1976 -101 1978 -99
rect 1980 -101 1981 -99
rect 1976 -106 1981 -101
rect 2004 -87 2012 -85
rect 2024 -86 2028 -77
rect 2004 -89 2005 -87
rect 2007 -89 2012 -87
rect 2004 -91 2012 -89
rect 2022 -87 2037 -86
rect 2022 -89 2024 -87
rect 2026 -89 2031 -87
rect 2033 -89 2037 -87
rect 2022 -90 2037 -89
rect 2007 -94 2012 -91
rect 2057 -87 2061 -74
rect 2057 -89 2058 -87
rect 2060 -89 2061 -87
rect 2007 -95 2045 -94
rect 2007 -97 2018 -95
rect 2020 -97 2045 -95
rect 2007 -98 2045 -97
rect 2057 -94 2061 -89
rect 2055 -96 2061 -94
rect 2055 -98 2056 -96
rect 2058 -98 2061 -96
rect 2055 -103 2061 -98
rect 2055 -105 2056 -103
rect 2058 -105 2061 -103
rect 1976 -108 1978 -106
rect 1980 -108 1981 -106
rect 1976 -110 1981 -108
rect 2055 -107 2061 -105
rect 2065 -71 2071 -70
rect 2065 -73 2068 -71
rect 2070 -73 2071 -71
rect 2065 -74 2071 -73
rect 2145 -70 2152 -69
rect 2145 -71 2149 -70
rect 2145 -73 2146 -71
rect 2148 -72 2149 -71
rect 2151 -72 2152 -70
rect 2148 -73 2152 -72
rect 2065 -94 2069 -74
rect 2098 -79 2102 -77
rect 2098 -81 2099 -79
rect 2101 -81 2102 -79
rect 2065 -96 2071 -94
rect 2065 -98 2068 -96
rect 2070 -98 2071 -96
rect 2065 -100 2071 -98
rect 2065 -102 2068 -100
rect 2070 -102 2071 -100
rect 2065 -103 2071 -102
rect 2065 -105 2068 -103
rect 2070 -105 2071 -103
rect 2065 -107 2071 -105
rect 2098 -86 2102 -81
rect 2145 -75 2150 -73
rect 2089 -87 2104 -86
rect 2089 -89 2093 -87
rect 2095 -89 2100 -87
rect 2102 -89 2104 -87
rect 2089 -90 2104 -89
rect 2114 -87 2122 -85
rect 2114 -89 2119 -87
rect 2121 -89 2122 -87
rect 2114 -91 2122 -89
rect 2114 -92 2119 -91
rect 2114 -94 2116 -92
rect 2118 -94 2119 -92
rect 2081 -98 2119 -94
rect 2146 -97 2150 -75
rect 2155 -81 2159 -77
rect 2155 -83 2156 -81
rect 2158 -83 2159 -81
rect 2155 -86 2159 -83
rect 2155 -87 2176 -86
rect 2155 -89 2170 -87
rect 2172 -89 2176 -87
rect 2155 -90 2176 -89
rect 2186 -78 2191 -76
rect 2186 -80 2187 -78
rect 2189 -80 2191 -78
rect 2186 -82 2191 -80
rect 2145 -99 2150 -97
rect 2145 -101 2146 -99
rect 2148 -101 2150 -99
rect 2145 -106 2150 -101
rect 2145 -108 2146 -106
rect 2148 -108 2150 -106
rect 2155 -96 2160 -94
rect 2162 -96 2176 -94
rect 2155 -98 2176 -96
rect 2155 -100 2159 -98
rect 2155 -102 2156 -100
rect 2158 -102 2159 -100
rect 2155 -107 2159 -102
rect 2145 -110 2150 -108
rect 2187 -101 2191 -82
rect 2255 -71 2259 -69
rect 2254 -73 2259 -71
rect 2254 -75 2255 -73
rect 2257 -75 2259 -73
rect 2254 -77 2259 -75
rect 2206 -79 2219 -78
rect 2206 -81 2210 -79
rect 2212 -81 2219 -79
rect 2206 -82 2219 -81
rect 2213 -87 2219 -82
rect 2213 -89 2214 -87
rect 2216 -89 2219 -87
rect 2213 -91 2219 -89
rect 2239 -92 2243 -85
rect 2239 -93 2241 -92
rect 2231 -94 2241 -93
rect 2231 -96 2236 -94
rect 2238 -96 2243 -94
rect 2231 -99 2243 -96
rect 2189 -103 2191 -101
rect 2187 -108 2191 -103
rect 2189 -110 2191 -108
rect 2178 -111 2191 -110
rect 2178 -113 2180 -111
rect 2182 -113 2191 -111
rect 2178 -114 2191 -113
rect 2187 -115 2191 -114
rect 2199 -106 2212 -102
rect 2199 -107 2204 -106
rect 2199 -109 2201 -107
rect 2203 -109 2204 -107
rect 2199 -115 2204 -109
rect 2255 -110 2259 -77
rect 2323 -71 2327 -69
rect 2322 -73 2327 -71
rect 2322 -75 2323 -73
rect 2325 -75 2327 -73
rect 2322 -77 2327 -75
rect 2274 -79 2287 -78
rect 2274 -81 2276 -79
rect 2278 -81 2287 -79
rect 2274 -82 2287 -81
rect 2281 -87 2287 -82
rect 2281 -89 2282 -87
rect 2284 -89 2287 -87
rect 2281 -91 2287 -89
rect 2307 -92 2311 -85
rect 2307 -93 2309 -92
rect 2299 -94 2309 -93
rect 2299 -96 2300 -94
rect 2302 -96 2311 -94
rect 2299 -99 2311 -96
rect 2246 -111 2259 -110
rect 2246 -113 2255 -111
rect 2257 -113 2259 -111
rect 2246 -114 2259 -113
rect 2267 -106 2280 -102
rect 2267 -107 2272 -106
rect 2267 -109 2269 -107
rect 2271 -109 2272 -107
rect 2267 -115 2272 -109
rect 2323 -110 2327 -77
rect 2314 -111 2327 -110
rect 2314 -113 2323 -111
rect 2325 -113 2327 -111
rect 2314 -114 2327 -113
rect 4 -121 2331 -120
rect 4 -123 39 -121
rect 41 -123 79 -121
rect 81 -123 298 -121
rect 300 -123 346 -121
rect 348 -123 565 -121
rect 567 -123 613 -121
rect 615 -123 832 -121
rect 834 -123 880 -121
rect 882 -123 1099 -121
rect 1101 -123 1147 -121
rect 1149 -123 1366 -121
rect 1368 -123 1414 -121
rect 1416 -123 1633 -121
rect 1635 -123 1681 -121
rect 1683 -123 1900 -121
rect 1902 -123 1948 -121
rect 1950 -123 2186 -121
rect 2188 -123 2320 -121
rect 2322 -123 2331 -121
rect 4 -133 2331 -123
rect 4 -135 39 -133
rect 41 -135 79 -133
rect 81 -135 298 -133
rect 300 -135 346 -133
rect 348 -135 565 -133
rect 567 -135 613 -133
rect 615 -135 832 -133
rect 834 -135 880 -133
rect 882 -135 1099 -133
rect 1101 -135 1147 -133
rect 1149 -135 1366 -133
rect 1368 -135 1414 -133
rect 1416 -135 1633 -133
rect 1635 -135 1681 -133
rect 1683 -135 1900 -133
rect 1902 -135 1948 -133
rect 1950 -135 2186 -133
rect 2188 -135 2331 -133
rect 4 -136 2331 -135
rect 8 -156 12 -149
rect 39 -147 44 -145
rect 39 -149 40 -147
rect 42 -149 44 -147
rect 8 -158 9 -156
rect 11 -158 12 -156
rect 8 -159 21 -158
rect 8 -161 13 -159
rect 15 -161 21 -159
rect 8 -162 21 -161
rect 15 -167 29 -166
rect 15 -169 23 -167
rect 25 -169 29 -167
rect 15 -170 29 -169
rect 39 -155 44 -149
rect 39 -157 40 -155
rect 42 -157 44 -155
rect 39 -159 44 -157
rect 39 -161 41 -159
rect 43 -161 44 -159
rect 39 -163 44 -161
rect 48 -158 52 -149
rect 299 -142 303 -141
rect 290 -146 303 -142
rect 88 -148 93 -146
rect 79 -150 84 -148
rect 48 -159 61 -158
rect 48 -161 53 -159
rect 55 -161 61 -159
rect 48 -162 61 -161
rect 15 -179 20 -170
rect 40 -181 44 -163
rect 55 -167 69 -166
rect 55 -169 63 -167
rect 65 -169 69 -167
rect 55 -170 69 -169
rect 79 -152 80 -150
rect 82 -152 84 -150
rect 79 -157 84 -152
rect 79 -159 80 -157
rect 82 -159 84 -157
rect 79 -161 84 -159
rect 55 -172 60 -170
rect 55 -174 57 -172
rect 59 -174 60 -172
rect 55 -179 60 -174
rect 80 -167 84 -161
rect 80 -169 81 -167
rect 83 -169 84 -167
rect 32 -183 40 -181
rect 42 -183 44 -181
rect 80 -181 84 -169
rect 32 -187 44 -183
rect 72 -183 80 -181
rect 82 -183 84 -181
rect 72 -187 84 -183
rect 88 -150 90 -148
rect 92 -150 93 -148
rect 88 -155 93 -150
rect 88 -157 90 -155
rect 92 -157 93 -155
rect 88 -159 93 -157
rect 88 -175 92 -159
rect 119 -159 157 -158
rect 119 -161 138 -159
rect 140 -161 157 -159
rect 119 -162 157 -161
rect 119 -165 124 -162
rect 116 -167 124 -165
rect 116 -169 117 -167
rect 119 -169 124 -167
rect 116 -171 124 -169
rect 134 -167 149 -166
rect 134 -169 136 -167
rect 138 -169 140 -167
rect 142 -169 143 -167
rect 145 -169 149 -167
rect 134 -170 149 -169
rect 88 -177 89 -175
rect 91 -177 92 -175
rect 88 -181 92 -177
rect 88 -183 93 -181
rect 136 -179 140 -170
rect 167 -151 173 -149
rect 167 -153 168 -151
rect 170 -153 173 -151
rect 167 -158 173 -153
rect 167 -160 168 -158
rect 170 -160 173 -158
rect 167 -162 173 -160
rect 169 -167 173 -162
rect 169 -169 170 -167
rect 172 -169 173 -167
rect 169 -182 173 -169
rect 88 -185 90 -183
rect 92 -185 93 -183
rect 88 -187 93 -185
rect 167 -183 173 -182
rect 167 -185 168 -183
rect 170 -185 173 -183
rect 167 -186 173 -185
rect 177 -151 183 -149
rect 257 -148 262 -146
rect 257 -150 258 -148
rect 260 -150 262 -148
rect 177 -153 180 -151
rect 182 -153 183 -151
rect 177 -154 183 -153
rect 177 -156 180 -154
rect 182 -156 183 -154
rect 177 -158 183 -156
rect 177 -160 180 -158
rect 182 -160 183 -158
rect 177 -162 183 -160
rect 177 -182 181 -162
rect 193 -159 231 -158
rect 193 -161 228 -159
rect 230 -161 231 -159
rect 193 -162 231 -161
rect 226 -165 231 -162
rect 201 -167 216 -166
rect 201 -169 205 -167
rect 207 -169 212 -167
rect 214 -169 216 -167
rect 201 -170 216 -169
rect 226 -167 234 -165
rect 226 -169 231 -167
rect 233 -169 234 -167
rect 210 -175 214 -170
rect 226 -171 234 -169
rect 257 -155 262 -150
rect 257 -157 258 -155
rect 260 -157 262 -155
rect 257 -159 262 -157
rect 210 -177 211 -175
rect 213 -177 214 -175
rect 210 -179 214 -177
rect 177 -183 183 -182
rect 177 -185 180 -183
rect 182 -185 183 -183
rect 177 -186 183 -185
rect 258 -181 262 -159
rect 267 -150 271 -149
rect 267 -152 268 -150
rect 270 -152 271 -150
rect 267 -158 271 -152
rect 267 -160 288 -158
rect 267 -162 272 -160
rect 274 -162 288 -160
rect 267 -167 288 -166
rect 267 -169 268 -167
rect 270 -169 282 -167
rect 284 -169 288 -167
rect 267 -170 288 -169
rect 301 -148 303 -146
rect 299 -153 303 -148
rect 301 -155 303 -153
rect 267 -174 271 -170
rect 299 -171 303 -155
rect 315 -158 319 -149
rect 566 -142 570 -141
rect 557 -146 570 -142
rect 355 -148 360 -146
rect 346 -150 351 -148
rect 315 -159 328 -158
rect 315 -161 320 -159
rect 322 -161 328 -159
rect 315 -162 328 -161
rect 299 -173 300 -171
rect 302 -173 303 -171
rect 299 -174 303 -173
rect 298 -176 303 -174
rect 298 -178 299 -176
rect 301 -178 303 -176
rect 298 -180 303 -178
rect 322 -167 336 -166
rect 322 -169 330 -167
rect 332 -169 336 -167
rect 322 -170 336 -169
rect 346 -152 347 -150
rect 349 -152 351 -150
rect 346 -157 351 -152
rect 346 -159 347 -157
rect 349 -159 351 -157
rect 346 -161 351 -159
rect 322 -172 327 -170
rect 322 -174 324 -172
rect 326 -174 327 -172
rect 322 -179 327 -174
rect 347 -167 351 -161
rect 347 -169 348 -167
rect 350 -169 351 -167
rect 257 -183 264 -181
rect 347 -181 351 -169
rect 257 -185 258 -183
rect 260 -184 264 -183
rect 260 -185 261 -184
rect 257 -186 261 -185
rect 263 -186 264 -184
rect 339 -183 347 -181
rect 349 -183 351 -181
rect 257 -187 264 -186
rect 339 -187 351 -183
rect 355 -150 357 -148
rect 359 -150 360 -148
rect 355 -155 360 -150
rect 355 -157 357 -155
rect 359 -157 360 -155
rect 355 -159 360 -157
rect 355 -175 359 -159
rect 386 -159 424 -158
rect 386 -161 405 -159
rect 407 -161 424 -159
rect 386 -162 424 -161
rect 386 -165 391 -162
rect 383 -167 391 -165
rect 383 -169 384 -167
rect 386 -169 391 -167
rect 383 -171 391 -169
rect 401 -167 416 -166
rect 401 -169 403 -167
rect 405 -169 407 -167
rect 409 -169 410 -167
rect 412 -169 416 -167
rect 401 -170 416 -169
rect 355 -177 356 -175
rect 358 -177 359 -175
rect 355 -181 359 -177
rect 355 -183 360 -181
rect 403 -179 407 -170
rect 434 -151 440 -149
rect 434 -153 435 -151
rect 437 -153 440 -151
rect 434 -158 440 -153
rect 434 -160 435 -158
rect 437 -160 440 -158
rect 434 -162 440 -160
rect 436 -167 440 -162
rect 436 -169 437 -167
rect 439 -169 440 -167
rect 436 -182 440 -169
rect 355 -185 357 -183
rect 359 -185 360 -183
rect 355 -187 360 -185
rect 434 -183 440 -182
rect 434 -185 435 -183
rect 437 -185 440 -183
rect 434 -186 440 -185
rect 444 -151 450 -149
rect 524 -148 529 -146
rect 524 -150 525 -148
rect 527 -150 529 -148
rect 444 -153 447 -151
rect 449 -153 450 -151
rect 444 -154 450 -153
rect 444 -156 447 -154
rect 449 -156 450 -154
rect 444 -158 450 -156
rect 444 -160 447 -158
rect 449 -160 450 -158
rect 444 -162 450 -160
rect 444 -182 448 -162
rect 460 -159 498 -158
rect 460 -161 495 -159
rect 497 -161 498 -159
rect 460 -162 498 -161
rect 493 -165 498 -162
rect 468 -167 483 -166
rect 468 -169 472 -167
rect 474 -169 479 -167
rect 481 -169 483 -167
rect 468 -170 483 -169
rect 493 -167 501 -165
rect 493 -169 498 -167
rect 500 -169 501 -167
rect 477 -175 481 -170
rect 493 -171 501 -169
rect 524 -155 529 -150
rect 524 -157 525 -155
rect 527 -157 529 -155
rect 524 -159 529 -157
rect 477 -177 478 -175
rect 480 -177 481 -175
rect 477 -179 481 -177
rect 444 -183 450 -182
rect 444 -185 447 -183
rect 449 -185 450 -183
rect 444 -186 450 -185
rect 525 -181 529 -159
rect 534 -150 538 -149
rect 534 -152 535 -150
rect 537 -152 538 -150
rect 534 -158 538 -152
rect 534 -160 555 -158
rect 534 -162 539 -160
rect 541 -162 555 -160
rect 534 -167 555 -166
rect 534 -169 535 -167
rect 537 -169 549 -167
rect 551 -169 555 -167
rect 534 -170 555 -169
rect 568 -148 570 -146
rect 566 -153 570 -148
rect 568 -155 570 -153
rect 534 -174 538 -170
rect 566 -171 570 -155
rect 582 -158 586 -149
rect 833 -142 837 -141
rect 824 -146 837 -142
rect 622 -148 627 -146
rect 613 -150 618 -148
rect 582 -159 595 -158
rect 582 -161 587 -159
rect 589 -161 595 -159
rect 582 -162 595 -161
rect 566 -173 567 -171
rect 569 -173 570 -171
rect 566 -174 570 -173
rect 565 -176 570 -174
rect 565 -178 566 -176
rect 568 -178 570 -176
rect 565 -180 570 -178
rect 589 -167 603 -166
rect 589 -169 597 -167
rect 599 -169 603 -167
rect 589 -170 603 -169
rect 613 -152 614 -150
rect 616 -152 618 -150
rect 613 -157 618 -152
rect 613 -159 614 -157
rect 616 -159 618 -157
rect 613 -161 618 -159
rect 589 -172 594 -170
rect 589 -174 591 -172
rect 593 -174 594 -172
rect 589 -179 594 -174
rect 614 -167 618 -161
rect 614 -169 615 -167
rect 617 -169 618 -167
rect 524 -183 531 -181
rect 614 -181 618 -169
rect 524 -185 525 -183
rect 527 -184 531 -183
rect 527 -185 528 -184
rect 524 -186 528 -185
rect 530 -186 531 -184
rect 606 -183 614 -181
rect 616 -183 618 -181
rect 524 -187 531 -186
rect 606 -187 618 -183
rect 622 -150 624 -148
rect 626 -150 627 -148
rect 622 -155 627 -150
rect 622 -157 624 -155
rect 626 -157 627 -155
rect 622 -159 627 -157
rect 622 -175 626 -159
rect 653 -159 691 -158
rect 653 -161 672 -159
rect 674 -161 691 -159
rect 653 -162 691 -161
rect 653 -165 658 -162
rect 650 -167 658 -165
rect 650 -169 651 -167
rect 653 -169 658 -167
rect 650 -171 658 -169
rect 668 -167 683 -166
rect 668 -169 670 -167
rect 672 -169 674 -167
rect 676 -169 677 -167
rect 679 -169 683 -167
rect 668 -170 683 -169
rect 622 -177 623 -175
rect 625 -177 626 -175
rect 622 -181 626 -177
rect 622 -183 627 -181
rect 670 -179 674 -170
rect 701 -151 707 -149
rect 701 -153 702 -151
rect 704 -153 707 -151
rect 701 -158 707 -153
rect 701 -160 702 -158
rect 704 -160 707 -158
rect 701 -162 707 -160
rect 703 -167 707 -162
rect 703 -169 704 -167
rect 706 -169 707 -167
rect 703 -182 707 -169
rect 622 -185 624 -183
rect 626 -185 627 -183
rect 622 -187 627 -185
rect 701 -183 707 -182
rect 701 -185 702 -183
rect 704 -185 707 -183
rect 701 -186 707 -185
rect 711 -151 717 -149
rect 791 -148 796 -146
rect 791 -150 792 -148
rect 794 -150 796 -148
rect 711 -153 714 -151
rect 716 -153 717 -151
rect 711 -154 717 -153
rect 711 -156 714 -154
rect 716 -156 717 -154
rect 711 -158 717 -156
rect 711 -160 714 -158
rect 716 -160 717 -158
rect 711 -162 717 -160
rect 711 -182 715 -162
rect 727 -159 765 -158
rect 727 -161 762 -159
rect 764 -161 765 -159
rect 727 -162 765 -161
rect 760 -165 765 -162
rect 735 -167 750 -166
rect 735 -169 739 -167
rect 741 -169 746 -167
rect 748 -169 750 -167
rect 735 -170 750 -169
rect 760 -167 768 -165
rect 760 -169 765 -167
rect 767 -169 768 -167
rect 744 -175 748 -170
rect 760 -171 768 -169
rect 791 -155 796 -150
rect 791 -157 792 -155
rect 794 -157 796 -155
rect 791 -159 796 -157
rect 744 -177 745 -175
rect 747 -177 748 -175
rect 744 -179 748 -177
rect 711 -183 717 -182
rect 711 -185 714 -183
rect 716 -185 717 -183
rect 711 -186 717 -185
rect 792 -181 796 -159
rect 801 -150 805 -149
rect 801 -152 802 -150
rect 804 -152 805 -150
rect 801 -158 805 -152
rect 801 -160 822 -158
rect 801 -162 806 -160
rect 808 -162 822 -160
rect 801 -167 822 -166
rect 801 -169 802 -167
rect 804 -169 816 -167
rect 818 -169 822 -167
rect 801 -170 822 -169
rect 835 -148 837 -146
rect 833 -153 837 -148
rect 835 -155 837 -153
rect 801 -174 805 -170
rect 833 -171 837 -155
rect 849 -158 853 -149
rect 1100 -142 1104 -141
rect 1091 -146 1104 -142
rect 889 -148 894 -146
rect 880 -150 885 -148
rect 849 -159 862 -158
rect 849 -161 854 -159
rect 856 -161 862 -159
rect 849 -162 862 -161
rect 833 -173 834 -171
rect 836 -173 837 -171
rect 833 -174 837 -173
rect 832 -176 837 -174
rect 832 -178 833 -176
rect 835 -178 837 -176
rect 832 -180 837 -178
rect 856 -167 870 -166
rect 856 -169 864 -167
rect 866 -169 870 -167
rect 856 -170 870 -169
rect 880 -152 881 -150
rect 883 -152 885 -150
rect 880 -157 885 -152
rect 880 -159 881 -157
rect 883 -159 885 -157
rect 880 -161 885 -159
rect 856 -172 861 -170
rect 856 -174 858 -172
rect 860 -174 861 -172
rect 856 -179 861 -174
rect 881 -167 885 -161
rect 881 -169 882 -167
rect 884 -169 885 -167
rect 791 -183 798 -181
rect 881 -181 885 -169
rect 791 -185 792 -183
rect 794 -184 798 -183
rect 794 -185 795 -184
rect 791 -186 795 -185
rect 797 -186 798 -184
rect 873 -183 881 -181
rect 883 -183 885 -181
rect 791 -187 798 -186
rect 873 -187 885 -183
rect 889 -150 891 -148
rect 893 -150 894 -148
rect 889 -155 894 -150
rect 889 -157 891 -155
rect 893 -157 894 -155
rect 889 -159 894 -157
rect 889 -175 893 -159
rect 920 -159 958 -158
rect 920 -161 939 -159
rect 941 -161 958 -159
rect 920 -162 958 -161
rect 920 -165 925 -162
rect 917 -167 925 -165
rect 917 -169 918 -167
rect 920 -169 925 -167
rect 917 -171 925 -169
rect 935 -167 950 -166
rect 935 -169 937 -167
rect 939 -169 941 -167
rect 943 -169 944 -167
rect 946 -169 950 -167
rect 935 -170 950 -169
rect 889 -177 890 -175
rect 892 -177 893 -175
rect 889 -181 893 -177
rect 889 -183 894 -181
rect 937 -179 941 -170
rect 968 -151 974 -149
rect 968 -153 969 -151
rect 971 -153 974 -151
rect 968 -158 974 -153
rect 968 -160 969 -158
rect 971 -160 974 -158
rect 968 -162 974 -160
rect 970 -167 974 -162
rect 970 -169 971 -167
rect 973 -169 974 -167
rect 970 -182 974 -169
rect 889 -185 891 -183
rect 893 -185 894 -183
rect 889 -187 894 -185
rect 968 -183 974 -182
rect 968 -185 969 -183
rect 971 -185 974 -183
rect 968 -186 974 -185
rect 978 -151 984 -149
rect 1058 -148 1063 -146
rect 1058 -150 1059 -148
rect 1061 -150 1063 -148
rect 978 -153 981 -151
rect 983 -153 984 -151
rect 978 -154 984 -153
rect 978 -156 981 -154
rect 983 -156 984 -154
rect 978 -158 984 -156
rect 978 -160 981 -158
rect 983 -160 984 -158
rect 978 -162 984 -160
rect 978 -182 982 -162
rect 994 -159 1032 -158
rect 994 -161 1029 -159
rect 1031 -161 1032 -159
rect 994 -162 1032 -161
rect 1027 -165 1032 -162
rect 1002 -167 1017 -166
rect 1002 -169 1006 -167
rect 1008 -169 1013 -167
rect 1015 -169 1017 -167
rect 1002 -170 1017 -169
rect 1027 -167 1035 -165
rect 1027 -169 1032 -167
rect 1034 -169 1035 -167
rect 1011 -175 1015 -170
rect 1027 -171 1035 -169
rect 1058 -155 1063 -150
rect 1058 -157 1059 -155
rect 1061 -157 1063 -155
rect 1058 -159 1063 -157
rect 1011 -177 1012 -175
rect 1014 -177 1015 -175
rect 1011 -179 1015 -177
rect 978 -183 984 -182
rect 978 -185 981 -183
rect 983 -185 984 -183
rect 978 -186 984 -185
rect 1059 -181 1063 -159
rect 1068 -150 1072 -149
rect 1068 -152 1069 -150
rect 1071 -152 1072 -150
rect 1068 -158 1072 -152
rect 1068 -160 1089 -158
rect 1068 -162 1073 -160
rect 1075 -162 1089 -160
rect 1068 -167 1089 -166
rect 1068 -169 1069 -167
rect 1071 -169 1083 -167
rect 1085 -169 1089 -167
rect 1068 -170 1089 -169
rect 1102 -148 1104 -146
rect 1100 -153 1104 -148
rect 1102 -155 1104 -153
rect 1068 -174 1072 -170
rect 1100 -171 1104 -155
rect 1116 -158 1120 -149
rect 1367 -142 1371 -141
rect 1358 -146 1371 -142
rect 1156 -148 1161 -146
rect 1147 -150 1152 -148
rect 1116 -159 1129 -158
rect 1116 -161 1121 -159
rect 1123 -161 1129 -159
rect 1116 -162 1129 -161
rect 1100 -173 1101 -171
rect 1103 -173 1104 -171
rect 1100 -174 1104 -173
rect 1099 -176 1104 -174
rect 1099 -178 1100 -176
rect 1102 -178 1104 -176
rect 1099 -180 1104 -178
rect 1123 -167 1137 -166
rect 1123 -169 1131 -167
rect 1133 -169 1137 -167
rect 1123 -170 1137 -169
rect 1147 -152 1148 -150
rect 1150 -152 1152 -150
rect 1147 -157 1152 -152
rect 1147 -159 1148 -157
rect 1150 -159 1152 -157
rect 1147 -161 1152 -159
rect 1123 -172 1128 -170
rect 1123 -174 1125 -172
rect 1127 -174 1128 -172
rect 1123 -179 1128 -174
rect 1148 -167 1152 -161
rect 1148 -169 1149 -167
rect 1151 -169 1152 -167
rect 1058 -183 1065 -181
rect 1148 -181 1152 -169
rect 1058 -185 1059 -183
rect 1061 -184 1065 -183
rect 1061 -185 1062 -184
rect 1058 -186 1062 -185
rect 1064 -186 1065 -184
rect 1140 -183 1148 -181
rect 1150 -183 1152 -181
rect 1058 -187 1065 -186
rect 1140 -187 1152 -183
rect 1156 -150 1158 -148
rect 1160 -150 1161 -148
rect 1156 -155 1161 -150
rect 1156 -157 1158 -155
rect 1160 -157 1161 -155
rect 1156 -159 1161 -157
rect 1156 -175 1160 -159
rect 1187 -159 1225 -158
rect 1187 -161 1206 -159
rect 1208 -161 1225 -159
rect 1187 -162 1225 -161
rect 1187 -165 1192 -162
rect 1184 -167 1192 -165
rect 1184 -169 1185 -167
rect 1187 -169 1192 -167
rect 1184 -171 1192 -169
rect 1202 -167 1217 -166
rect 1202 -169 1204 -167
rect 1206 -169 1208 -167
rect 1210 -169 1211 -167
rect 1213 -169 1217 -167
rect 1202 -170 1217 -169
rect 1156 -177 1157 -175
rect 1159 -177 1160 -175
rect 1156 -181 1160 -177
rect 1156 -183 1161 -181
rect 1204 -179 1208 -170
rect 1235 -151 1241 -149
rect 1235 -153 1236 -151
rect 1238 -153 1241 -151
rect 1235 -158 1241 -153
rect 1235 -160 1236 -158
rect 1238 -160 1241 -158
rect 1235 -162 1241 -160
rect 1237 -167 1241 -162
rect 1237 -169 1238 -167
rect 1240 -169 1241 -167
rect 1237 -182 1241 -169
rect 1156 -185 1158 -183
rect 1160 -185 1161 -183
rect 1156 -187 1161 -185
rect 1235 -183 1241 -182
rect 1235 -185 1236 -183
rect 1238 -185 1241 -183
rect 1235 -186 1241 -185
rect 1245 -151 1251 -149
rect 1325 -148 1330 -146
rect 1325 -150 1326 -148
rect 1328 -150 1330 -148
rect 1245 -153 1248 -151
rect 1250 -153 1251 -151
rect 1245 -154 1251 -153
rect 1245 -156 1248 -154
rect 1250 -156 1251 -154
rect 1245 -158 1251 -156
rect 1245 -160 1248 -158
rect 1250 -160 1251 -158
rect 1245 -162 1251 -160
rect 1245 -182 1249 -162
rect 1261 -159 1299 -158
rect 1261 -161 1296 -159
rect 1298 -161 1299 -159
rect 1261 -162 1299 -161
rect 1294 -165 1299 -162
rect 1269 -167 1284 -166
rect 1269 -169 1273 -167
rect 1275 -169 1280 -167
rect 1282 -169 1284 -167
rect 1269 -170 1284 -169
rect 1294 -167 1302 -165
rect 1294 -169 1299 -167
rect 1301 -169 1302 -167
rect 1278 -175 1282 -170
rect 1294 -171 1302 -169
rect 1325 -155 1330 -150
rect 1325 -157 1326 -155
rect 1328 -157 1330 -155
rect 1325 -159 1330 -157
rect 1278 -177 1279 -175
rect 1281 -177 1282 -175
rect 1278 -179 1282 -177
rect 1245 -183 1251 -182
rect 1245 -185 1248 -183
rect 1250 -185 1251 -183
rect 1245 -186 1251 -185
rect 1326 -181 1330 -159
rect 1335 -150 1339 -149
rect 1335 -152 1336 -150
rect 1338 -152 1339 -150
rect 1335 -158 1339 -152
rect 1335 -160 1356 -158
rect 1335 -162 1340 -160
rect 1342 -162 1356 -160
rect 1335 -167 1356 -166
rect 1335 -169 1336 -167
rect 1338 -169 1350 -167
rect 1352 -169 1356 -167
rect 1335 -170 1356 -169
rect 1369 -148 1371 -146
rect 1367 -153 1371 -148
rect 1369 -155 1371 -153
rect 1335 -174 1339 -170
rect 1367 -171 1371 -155
rect 1383 -158 1387 -149
rect 1634 -142 1638 -141
rect 1625 -146 1638 -142
rect 1423 -148 1428 -146
rect 1414 -150 1419 -148
rect 1383 -159 1396 -158
rect 1383 -161 1388 -159
rect 1390 -161 1396 -159
rect 1383 -162 1396 -161
rect 1367 -173 1368 -171
rect 1370 -173 1371 -171
rect 1367 -174 1371 -173
rect 1366 -176 1371 -174
rect 1366 -178 1367 -176
rect 1369 -178 1371 -176
rect 1366 -180 1371 -178
rect 1390 -167 1404 -166
rect 1390 -169 1398 -167
rect 1400 -169 1404 -167
rect 1390 -170 1404 -169
rect 1414 -152 1415 -150
rect 1417 -152 1419 -150
rect 1414 -157 1419 -152
rect 1414 -159 1415 -157
rect 1417 -159 1419 -157
rect 1414 -161 1419 -159
rect 1390 -172 1395 -170
rect 1390 -174 1392 -172
rect 1394 -174 1395 -172
rect 1390 -179 1395 -174
rect 1415 -167 1419 -161
rect 1415 -169 1416 -167
rect 1418 -169 1419 -167
rect 1325 -183 1332 -181
rect 1415 -181 1419 -169
rect 1325 -185 1326 -183
rect 1328 -184 1332 -183
rect 1328 -185 1329 -184
rect 1325 -186 1329 -185
rect 1331 -186 1332 -184
rect 1407 -183 1415 -181
rect 1417 -183 1419 -181
rect 1325 -187 1332 -186
rect 1407 -187 1419 -183
rect 1423 -150 1425 -148
rect 1427 -150 1428 -148
rect 1423 -155 1428 -150
rect 1423 -157 1425 -155
rect 1427 -157 1428 -155
rect 1423 -159 1428 -157
rect 1423 -175 1427 -159
rect 1454 -159 1492 -158
rect 1454 -161 1473 -159
rect 1475 -161 1492 -159
rect 1454 -162 1492 -161
rect 1454 -165 1459 -162
rect 1451 -167 1459 -165
rect 1451 -169 1452 -167
rect 1454 -169 1459 -167
rect 1451 -171 1459 -169
rect 1469 -167 1484 -166
rect 1469 -169 1471 -167
rect 1473 -169 1475 -167
rect 1477 -169 1478 -167
rect 1480 -169 1484 -167
rect 1469 -170 1484 -169
rect 1423 -177 1424 -175
rect 1426 -177 1427 -175
rect 1423 -181 1427 -177
rect 1423 -183 1428 -181
rect 1471 -179 1475 -170
rect 1502 -151 1508 -149
rect 1502 -153 1503 -151
rect 1505 -153 1508 -151
rect 1502 -158 1508 -153
rect 1502 -160 1503 -158
rect 1505 -160 1508 -158
rect 1502 -162 1508 -160
rect 1504 -167 1508 -162
rect 1504 -169 1505 -167
rect 1507 -169 1508 -167
rect 1504 -182 1508 -169
rect 1423 -185 1425 -183
rect 1427 -185 1428 -183
rect 1423 -187 1428 -185
rect 1502 -183 1508 -182
rect 1502 -185 1503 -183
rect 1505 -185 1508 -183
rect 1502 -186 1508 -185
rect 1512 -151 1518 -149
rect 1592 -148 1597 -146
rect 1592 -150 1593 -148
rect 1595 -150 1597 -148
rect 1512 -153 1515 -151
rect 1517 -153 1518 -151
rect 1512 -154 1518 -153
rect 1512 -156 1515 -154
rect 1517 -156 1518 -154
rect 1512 -158 1518 -156
rect 1512 -160 1515 -158
rect 1517 -160 1518 -158
rect 1512 -162 1518 -160
rect 1512 -182 1516 -162
rect 1528 -159 1566 -158
rect 1528 -161 1563 -159
rect 1565 -161 1566 -159
rect 1528 -162 1566 -161
rect 1561 -165 1566 -162
rect 1536 -167 1551 -166
rect 1536 -169 1540 -167
rect 1542 -169 1547 -167
rect 1549 -169 1551 -167
rect 1536 -170 1551 -169
rect 1561 -167 1569 -165
rect 1561 -169 1566 -167
rect 1568 -169 1569 -167
rect 1545 -175 1549 -170
rect 1561 -171 1569 -169
rect 1592 -155 1597 -150
rect 1592 -157 1593 -155
rect 1595 -157 1597 -155
rect 1592 -159 1597 -157
rect 1545 -177 1546 -175
rect 1548 -177 1549 -175
rect 1545 -179 1549 -177
rect 1512 -183 1518 -182
rect 1512 -185 1515 -183
rect 1517 -185 1518 -183
rect 1512 -186 1518 -185
rect 1593 -181 1597 -159
rect 1602 -150 1606 -149
rect 1602 -152 1603 -150
rect 1605 -152 1606 -150
rect 1602 -158 1606 -152
rect 1602 -160 1623 -158
rect 1602 -162 1607 -160
rect 1609 -162 1623 -160
rect 1602 -167 1623 -166
rect 1602 -169 1603 -167
rect 1605 -169 1617 -167
rect 1619 -169 1623 -167
rect 1602 -170 1623 -169
rect 1636 -148 1638 -146
rect 1634 -153 1638 -148
rect 1636 -155 1638 -153
rect 1602 -174 1606 -170
rect 1634 -171 1638 -155
rect 1650 -158 1654 -149
rect 1901 -142 1905 -141
rect 1892 -146 1905 -142
rect 1690 -148 1695 -146
rect 1681 -150 1686 -148
rect 1650 -159 1663 -158
rect 1650 -161 1655 -159
rect 1657 -161 1663 -159
rect 1650 -162 1663 -161
rect 1634 -173 1635 -171
rect 1637 -173 1638 -171
rect 1634 -174 1638 -173
rect 1633 -176 1638 -174
rect 1633 -178 1634 -176
rect 1636 -178 1638 -176
rect 1633 -180 1638 -178
rect 1657 -167 1671 -166
rect 1657 -169 1665 -167
rect 1667 -169 1671 -167
rect 1657 -170 1671 -169
rect 1681 -152 1682 -150
rect 1684 -152 1686 -150
rect 1681 -157 1686 -152
rect 1681 -159 1682 -157
rect 1684 -159 1686 -157
rect 1681 -161 1686 -159
rect 1657 -172 1662 -170
rect 1657 -174 1659 -172
rect 1661 -174 1662 -172
rect 1657 -179 1662 -174
rect 1682 -167 1686 -161
rect 1682 -169 1683 -167
rect 1685 -169 1686 -167
rect 1592 -183 1599 -181
rect 1682 -181 1686 -169
rect 1592 -185 1593 -183
rect 1595 -184 1599 -183
rect 1595 -185 1596 -184
rect 1592 -186 1596 -185
rect 1598 -186 1599 -184
rect 1674 -183 1682 -181
rect 1684 -183 1686 -181
rect 1592 -187 1599 -186
rect 1674 -187 1686 -183
rect 1690 -150 1692 -148
rect 1694 -150 1695 -148
rect 1690 -155 1695 -150
rect 1690 -157 1692 -155
rect 1694 -157 1695 -155
rect 1690 -159 1695 -157
rect 1690 -175 1694 -159
rect 1721 -159 1759 -158
rect 1721 -161 1740 -159
rect 1742 -161 1759 -159
rect 1721 -162 1759 -161
rect 1721 -165 1726 -162
rect 1718 -167 1726 -165
rect 1718 -169 1719 -167
rect 1721 -169 1726 -167
rect 1718 -171 1726 -169
rect 1736 -167 1751 -166
rect 1736 -169 1738 -167
rect 1740 -169 1742 -167
rect 1744 -169 1745 -167
rect 1747 -169 1751 -167
rect 1736 -170 1751 -169
rect 1690 -177 1691 -175
rect 1693 -177 1694 -175
rect 1690 -181 1694 -177
rect 1690 -183 1695 -181
rect 1738 -179 1742 -170
rect 1769 -151 1775 -149
rect 1769 -153 1770 -151
rect 1772 -153 1775 -151
rect 1769 -158 1775 -153
rect 1769 -160 1770 -158
rect 1772 -160 1775 -158
rect 1769 -162 1775 -160
rect 1771 -167 1775 -162
rect 1771 -169 1772 -167
rect 1774 -169 1775 -167
rect 1771 -182 1775 -169
rect 1690 -185 1692 -183
rect 1694 -185 1695 -183
rect 1690 -187 1695 -185
rect 1769 -183 1775 -182
rect 1769 -185 1770 -183
rect 1772 -185 1775 -183
rect 1769 -186 1775 -185
rect 1779 -151 1785 -149
rect 1859 -148 1864 -146
rect 1859 -150 1860 -148
rect 1862 -150 1864 -148
rect 1779 -153 1782 -151
rect 1784 -153 1785 -151
rect 1779 -154 1785 -153
rect 1779 -156 1782 -154
rect 1784 -156 1785 -154
rect 1779 -158 1785 -156
rect 1779 -160 1782 -158
rect 1784 -160 1785 -158
rect 1779 -162 1785 -160
rect 1779 -182 1783 -162
rect 1795 -159 1833 -158
rect 1795 -161 1830 -159
rect 1832 -161 1833 -159
rect 1795 -162 1833 -161
rect 1828 -165 1833 -162
rect 1803 -167 1818 -166
rect 1803 -169 1807 -167
rect 1809 -169 1814 -167
rect 1816 -169 1818 -167
rect 1803 -170 1818 -169
rect 1828 -167 1836 -165
rect 1828 -169 1833 -167
rect 1835 -169 1836 -167
rect 1812 -175 1816 -170
rect 1828 -171 1836 -169
rect 1859 -155 1864 -150
rect 1859 -157 1860 -155
rect 1862 -157 1864 -155
rect 1859 -159 1864 -157
rect 1812 -177 1813 -175
rect 1815 -177 1816 -175
rect 1812 -179 1816 -177
rect 1779 -183 1785 -182
rect 1779 -185 1782 -183
rect 1784 -185 1785 -183
rect 1779 -186 1785 -185
rect 1860 -176 1864 -159
rect 1869 -150 1873 -149
rect 1869 -152 1870 -150
rect 1872 -152 1873 -150
rect 1869 -158 1873 -152
rect 1869 -160 1890 -158
rect 1869 -162 1874 -160
rect 1876 -162 1890 -160
rect 1869 -167 1890 -166
rect 1869 -169 1870 -167
rect 1872 -169 1884 -167
rect 1886 -169 1890 -167
rect 1869 -170 1890 -169
rect 1903 -148 1905 -146
rect 1901 -153 1905 -148
rect 1903 -155 1905 -153
rect 1869 -174 1873 -170
rect 1901 -171 1905 -155
rect 1912 -147 1924 -141
rect 1912 -159 1917 -147
rect 2187 -142 2191 -141
rect 2178 -146 2191 -142
rect 1976 -148 1981 -146
rect 1912 -161 1914 -159
rect 1916 -161 1917 -159
rect 1912 -163 1917 -161
rect 1901 -173 1902 -171
rect 1904 -173 1905 -171
rect 1901 -174 1905 -173
rect 1860 -178 1861 -176
rect 1863 -178 1864 -176
rect 1860 -181 1864 -178
rect 1900 -176 1905 -174
rect 1900 -178 1901 -176
rect 1903 -178 1905 -176
rect 1900 -180 1905 -178
rect 1928 -172 1933 -165
rect 1956 -150 1972 -149
rect 1956 -152 1958 -150
rect 1960 -152 1972 -150
rect 1956 -154 1972 -152
rect 1968 -159 1972 -154
rect 1968 -161 1969 -159
rect 1971 -161 1972 -159
rect 1928 -173 1930 -172
rect 1920 -174 1930 -173
rect 1932 -174 1933 -172
rect 1920 -176 1933 -174
rect 1920 -178 1925 -176
rect 1927 -178 1933 -176
rect 1920 -179 1933 -178
rect 1859 -183 1866 -181
rect 1968 -182 1972 -161
rect 1859 -185 1860 -183
rect 1862 -185 1866 -183
rect 1859 -187 1866 -185
rect 1948 -183 1972 -182
rect 1948 -185 1950 -183
rect 1952 -185 1972 -183
rect 1948 -186 1972 -185
rect 1976 -150 1978 -148
rect 1980 -150 1981 -148
rect 1976 -155 1981 -150
rect 1976 -157 1978 -155
rect 1980 -157 1981 -155
rect 1976 -159 1981 -157
rect 1976 -175 1980 -159
rect 2007 -159 2045 -158
rect 2007 -161 2018 -159
rect 2020 -161 2045 -159
rect 2007 -162 2045 -161
rect 2007 -165 2012 -162
rect 2004 -167 2012 -165
rect 2004 -169 2005 -167
rect 2007 -169 2012 -167
rect 2004 -171 2012 -169
rect 2022 -167 2037 -166
rect 2022 -169 2024 -167
rect 2026 -169 2031 -167
rect 2033 -169 2037 -167
rect 2022 -170 2037 -169
rect 1976 -177 1977 -175
rect 1979 -177 1980 -175
rect 1976 -181 1980 -177
rect 1976 -183 1981 -181
rect 2024 -179 2028 -170
rect 2055 -151 2061 -149
rect 2055 -153 2056 -151
rect 2058 -153 2061 -151
rect 2055 -158 2061 -153
rect 2055 -160 2056 -158
rect 2058 -160 2061 -158
rect 2055 -162 2061 -160
rect 2057 -167 2061 -162
rect 2057 -169 2058 -167
rect 2060 -169 2061 -167
rect 2057 -182 2061 -169
rect 1976 -185 1978 -183
rect 1980 -185 1981 -183
rect 1976 -187 1981 -185
rect 2055 -183 2061 -182
rect 2055 -185 2056 -183
rect 2058 -185 2061 -183
rect 2055 -186 2061 -185
rect 2065 -151 2071 -149
rect 2145 -148 2150 -146
rect 2145 -150 2146 -148
rect 2148 -150 2150 -148
rect 2065 -153 2068 -151
rect 2070 -153 2071 -151
rect 2065 -154 2071 -153
rect 2065 -156 2068 -154
rect 2070 -156 2071 -154
rect 2065 -158 2071 -156
rect 2065 -160 2068 -158
rect 2070 -160 2071 -158
rect 2065 -162 2071 -160
rect 2065 -182 2069 -162
rect 2081 -159 2119 -158
rect 2081 -161 2116 -159
rect 2118 -161 2119 -159
rect 2081 -162 2119 -161
rect 2114 -165 2119 -162
rect 2089 -167 2104 -166
rect 2089 -169 2093 -167
rect 2095 -169 2100 -167
rect 2102 -169 2104 -167
rect 2089 -170 2104 -169
rect 2114 -167 2122 -165
rect 2114 -169 2119 -167
rect 2121 -169 2122 -167
rect 2098 -175 2102 -170
rect 2114 -171 2122 -169
rect 2145 -155 2150 -150
rect 2145 -157 2146 -155
rect 2148 -157 2150 -155
rect 2145 -159 2150 -157
rect 2098 -177 2099 -175
rect 2101 -177 2102 -175
rect 2098 -179 2102 -177
rect 2065 -183 2071 -182
rect 2065 -185 2068 -183
rect 2070 -185 2071 -183
rect 2065 -186 2071 -185
rect 2146 -179 2150 -159
rect 2155 -150 2159 -149
rect 2155 -152 2156 -150
rect 2158 -152 2159 -150
rect 2155 -158 2159 -152
rect 2155 -160 2176 -158
rect 2155 -162 2160 -160
rect 2162 -162 2176 -160
rect 2155 -167 2176 -166
rect 2155 -169 2156 -167
rect 2158 -169 2170 -167
rect 2172 -169 2176 -167
rect 2155 -170 2176 -169
rect 2189 -148 2191 -146
rect 2187 -153 2191 -148
rect 2189 -155 2191 -153
rect 2199 -147 2204 -141
rect 2246 -143 2259 -142
rect 2246 -145 2255 -143
rect 2257 -145 2259 -143
rect 2199 -149 2201 -147
rect 2203 -149 2204 -147
rect 2246 -146 2259 -145
rect 2199 -150 2204 -149
rect 2199 -154 2212 -150
rect 2155 -179 2159 -170
rect 2187 -171 2191 -155
rect 2187 -173 2188 -171
rect 2190 -173 2191 -171
rect 2187 -174 2191 -173
rect 2186 -176 2191 -174
rect 2186 -178 2187 -176
rect 2189 -178 2191 -176
rect 2146 -181 2147 -179
rect 2149 -181 2150 -179
rect 2186 -180 2191 -178
rect 2145 -183 2150 -181
rect 2145 -185 2146 -183
rect 2148 -185 2150 -183
rect 2213 -167 2219 -165
rect 2213 -169 2214 -167
rect 2216 -169 2219 -167
rect 2213 -174 2219 -169
rect 2206 -175 2219 -174
rect 2206 -177 2210 -175
rect 2212 -177 2219 -175
rect 2231 -158 2243 -157
rect 2231 -160 2236 -158
rect 2238 -160 2243 -158
rect 2231 -162 2243 -160
rect 2231 -163 2241 -162
rect 2239 -164 2241 -163
rect 2239 -171 2243 -164
rect 2206 -178 2219 -177
rect 2255 -179 2259 -146
rect 2267 -147 2272 -141
rect 2314 -143 2327 -142
rect 2314 -145 2323 -143
rect 2325 -145 2327 -143
rect 2267 -149 2269 -147
rect 2271 -149 2272 -147
rect 2314 -146 2327 -145
rect 2267 -150 2272 -149
rect 2267 -154 2280 -150
rect 2254 -181 2259 -179
rect 2145 -187 2150 -185
rect 2254 -183 2255 -181
rect 2257 -183 2259 -181
rect 2254 -185 2259 -183
rect 2281 -167 2287 -165
rect 2281 -169 2282 -167
rect 2284 -169 2287 -167
rect 2281 -174 2287 -169
rect 2274 -175 2287 -174
rect 2274 -177 2276 -175
rect 2278 -177 2287 -175
rect 2299 -158 2311 -157
rect 2299 -160 2300 -158
rect 2302 -160 2311 -158
rect 2299 -162 2311 -160
rect 2299 -163 2309 -162
rect 2307 -164 2309 -163
rect 2307 -171 2311 -164
rect 2274 -178 2287 -177
rect 2323 -179 2327 -146
rect 2322 -181 2327 -179
rect 2255 -187 2259 -185
rect 2322 -183 2323 -181
rect 2325 -183 2327 -181
rect 2322 -185 2327 -183
rect 2323 -187 2327 -185
rect 4 -193 2331 -192
rect 4 -195 29 -193
rect 31 -195 39 -193
rect 41 -195 69 -193
rect 71 -195 79 -193
rect 81 -195 298 -193
rect 300 -195 336 -193
rect 338 -195 346 -193
rect 348 -195 565 -193
rect 567 -195 603 -193
rect 605 -195 613 -193
rect 615 -195 832 -193
rect 834 -195 870 -193
rect 872 -195 880 -193
rect 882 -195 1099 -193
rect 1101 -195 1137 -193
rect 1139 -195 1147 -193
rect 1149 -195 1366 -193
rect 1368 -195 1404 -193
rect 1406 -195 1414 -193
rect 1416 -195 1633 -193
rect 1635 -195 1671 -193
rect 1673 -195 1681 -193
rect 1683 -195 1900 -193
rect 1902 -195 1915 -193
rect 1917 -195 1968 -193
rect 1970 -195 2186 -193
rect 2188 -195 2324 -193
rect 2326 -195 2331 -193
rect 4 -199 2331 -195
rect 4 -201 2276 -199
rect 2278 -201 2331 -199
rect 4 -202 2331 -201
rect 4 -204 133 -202
rect 135 -204 400 -202
rect 402 -204 667 -202
rect 669 -204 934 -202
rect 936 -204 1201 -202
rect 1203 -204 1468 -202
rect 1470 -204 1735 -202
rect 1737 -204 2331 -202
rect 4 -205 2331 -204
rect 4 -207 29 -205
rect 31 -207 39 -205
rect 41 -207 69 -205
rect 71 -207 79 -205
rect 81 -207 298 -205
rect 300 -207 336 -205
rect 338 -207 346 -205
rect 348 -207 565 -205
rect 567 -207 603 -205
rect 605 -207 613 -205
rect 615 -207 832 -205
rect 834 -207 870 -205
rect 872 -207 880 -205
rect 882 -207 1099 -205
rect 1101 -207 1137 -205
rect 1139 -207 1147 -205
rect 1149 -207 1366 -205
rect 1368 -207 1404 -205
rect 1406 -207 1414 -205
rect 1416 -207 1633 -205
rect 1635 -207 1671 -205
rect 1673 -207 1681 -205
rect 1683 -207 1900 -205
rect 1902 -207 1915 -205
rect 1917 -207 1968 -205
rect 1970 -207 2186 -205
rect 2188 -207 2331 -205
rect 4 -208 2331 -207
rect 15 -230 20 -221
rect 32 -217 44 -213
rect 32 -219 40 -217
rect 42 -219 44 -217
rect 15 -231 29 -230
rect 15 -233 23 -231
rect 25 -233 29 -231
rect 15 -234 29 -233
rect 8 -239 21 -238
rect 8 -241 13 -239
rect 15 -241 21 -239
rect 8 -242 21 -241
rect 8 -243 12 -242
rect 8 -245 9 -243
rect 11 -245 12 -243
rect 40 -231 44 -219
rect 40 -233 41 -231
rect 43 -233 44 -231
rect 40 -239 44 -233
rect 55 -230 60 -221
rect 72 -217 84 -213
rect 72 -219 80 -217
rect 82 -219 84 -217
rect 55 -231 69 -230
rect 55 -233 63 -231
rect 65 -233 69 -231
rect 55 -234 69 -233
rect 8 -251 12 -245
rect 39 -241 44 -239
rect 39 -243 40 -241
rect 42 -243 44 -241
rect 39 -248 44 -243
rect 39 -250 40 -248
rect 42 -250 44 -248
rect 39 -252 44 -250
rect 48 -239 61 -238
rect 48 -241 53 -239
rect 55 -241 61 -239
rect 48 -242 61 -241
rect 48 -244 52 -242
rect 48 -246 49 -244
rect 51 -246 52 -244
rect 80 -231 84 -219
rect 80 -233 81 -231
rect 83 -233 84 -231
rect 80 -239 84 -233
rect 48 -251 52 -246
rect 79 -241 84 -239
rect 79 -243 80 -241
rect 82 -243 84 -241
rect 79 -248 84 -243
rect 79 -250 80 -248
rect 82 -250 84 -248
rect 79 -252 84 -250
rect 88 -215 93 -213
rect 88 -217 90 -215
rect 92 -217 93 -215
rect 88 -219 93 -217
rect 88 -223 92 -219
rect 88 -225 89 -223
rect 91 -225 92 -223
rect 88 -241 92 -225
rect 167 -215 173 -214
rect 167 -217 168 -215
rect 170 -217 173 -215
rect 167 -218 173 -217
rect 88 -243 93 -241
rect 88 -245 90 -243
rect 92 -245 93 -243
rect 88 -250 93 -245
rect 116 -231 124 -229
rect 136 -230 140 -221
rect 116 -233 117 -231
rect 119 -233 124 -231
rect 116 -235 124 -233
rect 134 -231 149 -230
rect 134 -233 136 -231
rect 138 -233 139 -231
rect 141 -233 143 -231
rect 145 -233 149 -231
rect 134 -234 149 -233
rect 119 -238 124 -235
rect 169 -231 173 -218
rect 169 -233 170 -231
rect 172 -233 173 -231
rect 119 -239 157 -238
rect 119 -241 133 -239
rect 135 -241 157 -239
rect 119 -242 157 -241
rect 169 -238 173 -233
rect 167 -240 173 -238
rect 167 -242 168 -240
rect 170 -242 173 -240
rect 167 -247 173 -242
rect 167 -249 168 -247
rect 170 -249 173 -247
rect 88 -252 90 -250
rect 92 -252 93 -250
rect 88 -254 93 -252
rect 167 -251 173 -249
rect 177 -215 183 -214
rect 177 -217 180 -215
rect 182 -217 183 -215
rect 177 -218 183 -217
rect 257 -214 264 -213
rect 257 -215 261 -214
rect 257 -217 258 -215
rect 260 -216 261 -215
rect 263 -216 264 -214
rect 260 -217 264 -216
rect 177 -238 181 -218
rect 210 -223 214 -221
rect 210 -225 211 -223
rect 213 -225 214 -223
rect 177 -240 183 -238
rect 177 -242 180 -240
rect 182 -242 183 -240
rect 177 -244 183 -242
rect 177 -246 180 -244
rect 182 -246 183 -244
rect 177 -247 183 -246
rect 177 -249 180 -247
rect 182 -249 183 -247
rect 177 -251 183 -249
rect 210 -230 214 -225
rect 257 -219 264 -217
rect 201 -231 216 -230
rect 201 -233 205 -231
rect 207 -233 212 -231
rect 214 -233 216 -231
rect 201 -234 216 -233
rect 226 -231 234 -229
rect 226 -233 231 -231
rect 233 -233 234 -231
rect 226 -235 234 -233
rect 226 -236 231 -235
rect 226 -238 228 -236
rect 230 -238 231 -236
rect 193 -242 231 -238
rect 258 -241 262 -219
rect 267 -225 271 -224
rect 267 -227 268 -225
rect 270 -227 271 -225
rect 267 -230 271 -227
rect 267 -231 288 -230
rect 267 -233 282 -231
rect 284 -233 288 -231
rect 267 -234 288 -233
rect 298 -222 303 -220
rect 298 -224 299 -222
rect 301 -224 303 -222
rect 298 -226 303 -224
rect 257 -243 262 -241
rect 257 -245 258 -243
rect 260 -245 262 -243
rect 257 -250 262 -245
rect 257 -252 258 -250
rect 260 -252 262 -250
rect 267 -240 272 -238
rect 274 -240 288 -238
rect 267 -242 288 -240
rect 267 -244 271 -242
rect 267 -246 268 -244
rect 270 -246 271 -244
rect 267 -251 271 -246
rect 257 -254 262 -252
rect 299 -245 303 -226
rect 322 -230 327 -221
rect 339 -217 351 -213
rect 339 -219 347 -217
rect 349 -219 351 -217
rect 322 -231 336 -230
rect 322 -233 330 -231
rect 332 -233 336 -231
rect 322 -234 336 -233
rect 301 -247 303 -245
rect 299 -252 303 -247
rect 315 -239 328 -238
rect 315 -241 320 -239
rect 322 -241 328 -239
rect 315 -242 328 -241
rect 315 -244 319 -242
rect 315 -246 316 -244
rect 318 -246 319 -244
rect 347 -231 351 -219
rect 347 -233 348 -231
rect 350 -233 351 -231
rect 347 -239 351 -233
rect 315 -251 319 -246
rect 346 -241 351 -239
rect 346 -243 347 -241
rect 349 -243 351 -241
rect 346 -248 351 -243
rect 301 -254 303 -252
rect 290 -256 303 -254
rect 290 -258 300 -256
rect 302 -258 303 -256
rect 299 -259 303 -258
rect 346 -250 347 -248
rect 349 -250 351 -248
rect 346 -252 351 -250
rect 355 -215 360 -213
rect 355 -217 357 -215
rect 359 -217 360 -215
rect 355 -219 360 -217
rect 355 -223 359 -219
rect 355 -225 356 -223
rect 358 -225 359 -223
rect 355 -241 359 -225
rect 434 -215 440 -214
rect 434 -217 435 -215
rect 437 -217 440 -215
rect 434 -218 440 -217
rect 355 -243 360 -241
rect 355 -245 357 -243
rect 359 -245 360 -243
rect 355 -250 360 -245
rect 383 -231 391 -229
rect 403 -230 407 -221
rect 383 -233 384 -231
rect 386 -233 391 -231
rect 383 -235 391 -233
rect 401 -231 416 -230
rect 401 -233 403 -231
rect 405 -233 406 -231
rect 408 -233 410 -231
rect 412 -233 416 -231
rect 401 -234 416 -233
rect 386 -238 391 -235
rect 436 -231 440 -218
rect 436 -233 437 -231
rect 439 -233 440 -231
rect 386 -239 424 -238
rect 386 -241 400 -239
rect 402 -241 424 -239
rect 386 -242 424 -241
rect 436 -238 440 -233
rect 434 -240 440 -238
rect 434 -242 435 -240
rect 437 -242 440 -240
rect 434 -247 440 -242
rect 434 -249 435 -247
rect 437 -249 440 -247
rect 355 -252 357 -250
rect 359 -252 360 -250
rect 355 -254 360 -252
rect 434 -251 440 -249
rect 444 -215 450 -214
rect 444 -217 447 -215
rect 449 -217 450 -215
rect 444 -218 450 -217
rect 524 -214 531 -213
rect 524 -215 528 -214
rect 524 -217 525 -215
rect 527 -216 528 -215
rect 530 -216 531 -214
rect 527 -217 531 -216
rect 444 -238 448 -218
rect 477 -223 481 -221
rect 477 -225 478 -223
rect 480 -225 481 -223
rect 444 -240 450 -238
rect 444 -242 447 -240
rect 449 -242 450 -240
rect 444 -244 450 -242
rect 444 -246 447 -244
rect 449 -246 450 -244
rect 444 -247 450 -246
rect 444 -249 447 -247
rect 449 -249 450 -247
rect 444 -251 450 -249
rect 477 -230 481 -225
rect 524 -219 531 -217
rect 468 -231 483 -230
rect 468 -233 472 -231
rect 474 -233 479 -231
rect 481 -233 483 -231
rect 468 -234 483 -233
rect 493 -231 501 -229
rect 493 -233 498 -231
rect 500 -233 501 -231
rect 493 -235 501 -233
rect 493 -236 498 -235
rect 493 -238 495 -236
rect 497 -238 498 -236
rect 460 -242 498 -238
rect 525 -241 529 -219
rect 534 -225 538 -224
rect 534 -227 535 -225
rect 537 -227 538 -225
rect 534 -230 538 -227
rect 534 -231 555 -230
rect 534 -233 549 -231
rect 551 -233 555 -231
rect 534 -234 555 -233
rect 565 -222 570 -220
rect 565 -224 566 -222
rect 568 -224 570 -222
rect 565 -226 570 -224
rect 524 -243 529 -241
rect 524 -245 525 -243
rect 527 -245 529 -243
rect 524 -250 529 -245
rect 524 -252 525 -250
rect 527 -252 529 -250
rect 534 -240 539 -238
rect 541 -240 555 -238
rect 534 -242 555 -240
rect 534 -244 538 -242
rect 534 -246 535 -244
rect 537 -246 538 -244
rect 534 -251 538 -246
rect 524 -254 529 -252
rect 566 -245 570 -226
rect 589 -230 594 -221
rect 606 -217 618 -213
rect 606 -219 614 -217
rect 616 -219 618 -217
rect 589 -231 603 -230
rect 589 -233 597 -231
rect 599 -233 603 -231
rect 589 -234 603 -233
rect 568 -247 570 -245
rect 566 -252 570 -247
rect 582 -239 595 -238
rect 582 -241 587 -239
rect 589 -241 595 -239
rect 582 -242 595 -241
rect 582 -244 586 -242
rect 582 -246 583 -244
rect 585 -246 586 -244
rect 614 -231 618 -219
rect 614 -233 615 -231
rect 617 -233 618 -231
rect 614 -239 618 -233
rect 582 -251 586 -246
rect 613 -241 618 -239
rect 613 -243 614 -241
rect 616 -243 618 -241
rect 613 -248 618 -243
rect 568 -254 570 -252
rect 557 -256 570 -254
rect 557 -258 567 -256
rect 569 -258 570 -256
rect 566 -259 570 -258
rect 613 -250 614 -248
rect 616 -250 618 -248
rect 613 -252 618 -250
rect 622 -215 627 -213
rect 622 -217 624 -215
rect 626 -217 627 -215
rect 622 -219 627 -217
rect 622 -223 626 -219
rect 622 -225 623 -223
rect 625 -225 626 -223
rect 622 -241 626 -225
rect 701 -215 707 -214
rect 701 -217 702 -215
rect 704 -217 707 -215
rect 701 -218 707 -217
rect 622 -243 627 -241
rect 622 -245 624 -243
rect 626 -245 627 -243
rect 622 -250 627 -245
rect 650 -231 658 -229
rect 670 -230 674 -221
rect 650 -233 651 -231
rect 653 -233 658 -231
rect 650 -235 658 -233
rect 668 -231 683 -230
rect 668 -233 670 -231
rect 672 -233 673 -231
rect 675 -233 677 -231
rect 679 -233 683 -231
rect 668 -234 683 -233
rect 653 -238 658 -235
rect 703 -231 707 -218
rect 703 -233 704 -231
rect 706 -233 707 -231
rect 653 -239 691 -238
rect 653 -241 667 -239
rect 669 -241 691 -239
rect 653 -242 691 -241
rect 703 -238 707 -233
rect 701 -240 707 -238
rect 701 -242 702 -240
rect 704 -242 707 -240
rect 701 -247 707 -242
rect 701 -249 702 -247
rect 704 -249 707 -247
rect 622 -252 624 -250
rect 626 -252 627 -250
rect 622 -254 627 -252
rect 701 -251 707 -249
rect 711 -215 717 -214
rect 711 -217 714 -215
rect 716 -217 717 -215
rect 711 -218 717 -217
rect 791 -214 798 -213
rect 791 -215 795 -214
rect 791 -217 792 -215
rect 794 -216 795 -215
rect 797 -216 798 -214
rect 794 -217 798 -216
rect 711 -238 715 -218
rect 744 -223 748 -221
rect 744 -225 745 -223
rect 747 -225 748 -223
rect 711 -240 717 -238
rect 711 -242 714 -240
rect 716 -242 717 -240
rect 711 -244 717 -242
rect 711 -246 714 -244
rect 716 -246 717 -244
rect 711 -247 717 -246
rect 711 -249 714 -247
rect 716 -249 717 -247
rect 711 -251 717 -249
rect 744 -230 748 -225
rect 791 -219 798 -217
rect 735 -231 750 -230
rect 735 -233 739 -231
rect 741 -233 746 -231
rect 748 -233 750 -231
rect 735 -234 750 -233
rect 760 -231 768 -229
rect 760 -233 765 -231
rect 767 -233 768 -231
rect 760 -235 768 -233
rect 760 -236 765 -235
rect 760 -238 762 -236
rect 764 -238 765 -236
rect 727 -242 765 -238
rect 792 -241 796 -219
rect 801 -225 805 -224
rect 801 -227 802 -225
rect 804 -227 805 -225
rect 801 -230 805 -227
rect 801 -231 822 -230
rect 801 -233 816 -231
rect 818 -233 822 -231
rect 801 -234 822 -233
rect 832 -222 837 -220
rect 832 -224 833 -222
rect 835 -224 837 -222
rect 832 -226 837 -224
rect 791 -243 796 -241
rect 791 -245 792 -243
rect 794 -245 796 -243
rect 791 -250 796 -245
rect 791 -252 792 -250
rect 794 -252 796 -250
rect 801 -240 806 -238
rect 808 -240 822 -238
rect 801 -242 822 -240
rect 801 -244 805 -242
rect 801 -246 802 -244
rect 804 -246 805 -244
rect 801 -251 805 -246
rect 791 -254 796 -252
rect 833 -245 837 -226
rect 856 -230 861 -221
rect 873 -217 885 -213
rect 873 -219 881 -217
rect 883 -219 885 -217
rect 856 -231 870 -230
rect 856 -233 864 -231
rect 866 -233 870 -231
rect 856 -234 870 -233
rect 835 -247 837 -245
rect 833 -252 837 -247
rect 849 -239 862 -238
rect 849 -241 854 -239
rect 856 -241 862 -239
rect 849 -242 862 -241
rect 849 -244 853 -242
rect 849 -246 850 -244
rect 852 -246 853 -244
rect 881 -231 885 -219
rect 881 -233 882 -231
rect 884 -233 885 -231
rect 881 -239 885 -233
rect 849 -251 853 -246
rect 880 -241 885 -239
rect 880 -243 881 -241
rect 883 -243 885 -241
rect 880 -248 885 -243
rect 835 -254 837 -252
rect 824 -256 837 -254
rect 824 -258 834 -256
rect 836 -258 837 -256
rect 833 -259 837 -258
rect 880 -250 881 -248
rect 883 -250 885 -248
rect 880 -252 885 -250
rect 889 -215 894 -213
rect 889 -217 891 -215
rect 893 -217 894 -215
rect 889 -219 894 -217
rect 889 -223 893 -219
rect 889 -225 890 -223
rect 892 -225 893 -223
rect 889 -241 893 -225
rect 968 -215 974 -214
rect 968 -217 969 -215
rect 971 -217 974 -215
rect 968 -218 974 -217
rect 889 -243 894 -241
rect 889 -245 891 -243
rect 893 -245 894 -243
rect 889 -250 894 -245
rect 917 -231 925 -229
rect 937 -230 941 -221
rect 917 -233 918 -231
rect 920 -233 925 -231
rect 917 -235 925 -233
rect 935 -231 950 -230
rect 935 -233 937 -231
rect 939 -233 940 -231
rect 942 -233 944 -231
rect 946 -233 950 -231
rect 935 -234 950 -233
rect 920 -238 925 -235
rect 970 -231 974 -218
rect 970 -233 971 -231
rect 973 -233 974 -231
rect 920 -239 958 -238
rect 920 -241 934 -239
rect 936 -241 958 -239
rect 920 -242 958 -241
rect 970 -238 974 -233
rect 968 -240 974 -238
rect 968 -242 969 -240
rect 971 -242 974 -240
rect 968 -247 974 -242
rect 968 -249 969 -247
rect 971 -249 974 -247
rect 889 -252 891 -250
rect 893 -252 894 -250
rect 889 -254 894 -252
rect 968 -251 974 -249
rect 978 -215 984 -214
rect 978 -217 981 -215
rect 983 -217 984 -215
rect 978 -218 984 -217
rect 1058 -214 1065 -213
rect 1058 -215 1062 -214
rect 1058 -217 1059 -215
rect 1061 -216 1062 -215
rect 1064 -216 1065 -214
rect 1061 -217 1065 -216
rect 978 -238 982 -218
rect 1011 -223 1015 -221
rect 1011 -225 1012 -223
rect 1014 -225 1015 -223
rect 978 -240 984 -238
rect 978 -242 981 -240
rect 983 -242 984 -240
rect 978 -244 984 -242
rect 978 -246 981 -244
rect 983 -246 984 -244
rect 978 -247 984 -246
rect 978 -249 981 -247
rect 983 -249 984 -247
rect 978 -251 984 -249
rect 1011 -230 1015 -225
rect 1058 -219 1065 -217
rect 1002 -231 1017 -230
rect 1002 -233 1006 -231
rect 1008 -233 1013 -231
rect 1015 -233 1017 -231
rect 1002 -234 1017 -233
rect 1027 -231 1035 -229
rect 1027 -233 1032 -231
rect 1034 -233 1035 -231
rect 1027 -235 1035 -233
rect 1027 -236 1032 -235
rect 1027 -238 1029 -236
rect 1031 -238 1032 -236
rect 994 -242 1032 -238
rect 1059 -241 1063 -219
rect 1068 -225 1072 -224
rect 1068 -227 1069 -225
rect 1071 -227 1072 -225
rect 1068 -230 1072 -227
rect 1068 -231 1089 -230
rect 1068 -233 1083 -231
rect 1085 -233 1089 -231
rect 1068 -234 1089 -233
rect 1099 -222 1104 -220
rect 1099 -224 1100 -222
rect 1102 -224 1104 -222
rect 1099 -226 1104 -224
rect 1058 -243 1063 -241
rect 1058 -245 1059 -243
rect 1061 -245 1063 -243
rect 1058 -250 1063 -245
rect 1058 -252 1059 -250
rect 1061 -252 1063 -250
rect 1068 -240 1073 -238
rect 1075 -240 1089 -238
rect 1068 -242 1089 -240
rect 1068 -244 1072 -242
rect 1068 -246 1069 -244
rect 1071 -246 1072 -244
rect 1068 -251 1072 -246
rect 1058 -254 1063 -252
rect 1100 -245 1104 -226
rect 1123 -230 1128 -221
rect 1140 -217 1152 -213
rect 1140 -219 1148 -217
rect 1150 -219 1152 -217
rect 1123 -231 1137 -230
rect 1123 -233 1131 -231
rect 1133 -233 1137 -231
rect 1123 -234 1137 -233
rect 1102 -247 1104 -245
rect 1100 -252 1104 -247
rect 1116 -239 1129 -238
rect 1116 -241 1121 -239
rect 1123 -241 1129 -239
rect 1116 -242 1129 -241
rect 1116 -244 1120 -242
rect 1116 -246 1117 -244
rect 1119 -246 1120 -244
rect 1148 -231 1152 -219
rect 1148 -233 1149 -231
rect 1151 -233 1152 -231
rect 1148 -239 1152 -233
rect 1116 -251 1120 -246
rect 1147 -241 1152 -239
rect 1147 -243 1148 -241
rect 1150 -243 1152 -241
rect 1147 -248 1152 -243
rect 1102 -254 1104 -252
rect 1091 -256 1104 -254
rect 1091 -258 1101 -256
rect 1103 -258 1104 -256
rect 1100 -259 1104 -258
rect 1147 -250 1148 -248
rect 1150 -250 1152 -248
rect 1147 -252 1152 -250
rect 1156 -215 1161 -213
rect 1156 -217 1158 -215
rect 1160 -217 1161 -215
rect 1156 -219 1161 -217
rect 1156 -223 1160 -219
rect 1156 -225 1157 -223
rect 1159 -225 1160 -223
rect 1156 -241 1160 -225
rect 1235 -215 1241 -214
rect 1235 -217 1236 -215
rect 1238 -217 1241 -215
rect 1235 -218 1241 -217
rect 1156 -243 1161 -241
rect 1156 -245 1158 -243
rect 1160 -245 1161 -243
rect 1156 -250 1161 -245
rect 1184 -231 1192 -229
rect 1204 -230 1208 -221
rect 1184 -233 1185 -231
rect 1187 -233 1192 -231
rect 1184 -235 1192 -233
rect 1202 -231 1217 -230
rect 1202 -233 1204 -231
rect 1206 -233 1207 -231
rect 1209 -233 1211 -231
rect 1213 -233 1217 -231
rect 1202 -234 1217 -233
rect 1187 -238 1192 -235
rect 1237 -231 1241 -218
rect 1237 -233 1238 -231
rect 1240 -233 1241 -231
rect 1187 -239 1225 -238
rect 1187 -241 1201 -239
rect 1203 -241 1225 -239
rect 1187 -242 1225 -241
rect 1237 -238 1241 -233
rect 1235 -240 1241 -238
rect 1235 -242 1236 -240
rect 1238 -242 1241 -240
rect 1235 -247 1241 -242
rect 1235 -249 1236 -247
rect 1238 -249 1241 -247
rect 1156 -252 1158 -250
rect 1160 -252 1161 -250
rect 1156 -254 1161 -252
rect 1235 -251 1241 -249
rect 1245 -215 1251 -214
rect 1245 -217 1248 -215
rect 1250 -217 1251 -215
rect 1245 -218 1251 -217
rect 1325 -214 1332 -213
rect 1325 -215 1329 -214
rect 1325 -217 1326 -215
rect 1328 -216 1329 -215
rect 1331 -216 1332 -214
rect 1328 -217 1332 -216
rect 1245 -238 1249 -218
rect 1278 -223 1282 -221
rect 1278 -225 1279 -223
rect 1281 -225 1282 -223
rect 1245 -240 1251 -238
rect 1245 -242 1248 -240
rect 1250 -242 1251 -240
rect 1245 -244 1251 -242
rect 1245 -246 1248 -244
rect 1250 -246 1251 -244
rect 1245 -247 1251 -246
rect 1245 -249 1248 -247
rect 1250 -249 1251 -247
rect 1245 -251 1251 -249
rect 1278 -230 1282 -225
rect 1325 -219 1332 -217
rect 1269 -231 1284 -230
rect 1269 -233 1273 -231
rect 1275 -233 1280 -231
rect 1282 -233 1284 -231
rect 1269 -234 1284 -233
rect 1294 -231 1302 -229
rect 1294 -233 1299 -231
rect 1301 -233 1302 -231
rect 1294 -235 1302 -233
rect 1294 -236 1299 -235
rect 1294 -238 1296 -236
rect 1298 -238 1299 -236
rect 1261 -242 1299 -238
rect 1326 -241 1330 -219
rect 1335 -225 1339 -224
rect 1335 -227 1336 -225
rect 1338 -227 1339 -225
rect 1335 -230 1339 -227
rect 1335 -231 1356 -230
rect 1335 -233 1350 -231
rect 1352 -233 1356 -231
rect 1335 -234 1356 -233
rect 1366 -222 1371 -220
rect 1366 -224 1367 -222
rect 1369 -224 1371 -222
rect 1366 -226 1371 -224
rect 1325 -243 1330 -241
rect 1325 -245 1326 -243
rect 1328 -245 1330 -243
rect 1325 -250 1330 -245
rect 1325 -252 1326 -250
rect 1328 -252 1330 -250
rect 1335 -240 1340 -238
rect 1342 -240 1356 -238
rect 1335 -242 1356 -240
rect 1335 -244 1339 -242
rect 1335 -246 1336 -244
rect 1338 -246 1339 -244
rect 1335 -251 1339 -246
rect 1325 -254 1330 -252
rect 1367 -245 1371 -226
rect 1390 -230 1395 -221
rect 1407 -217 1419 -213
rect 1407 -219 1415 -217
rect 1417 -219 1419 -217
rect 1390 -231 1404 -230
rect 1390 -233 1398 -231
rect 1400 -233 1404 -231
rect 1390 -234 1404 -233
rect 1369 -247 1371 -245
rect 1367 -252 1371 -247
rect 1383 -239 1396 -238
rect 1383 -241 1388 -239
rect 1390 -241 1396 -239
rect 1383 -242 1396 -241
rect 1383 -244 1387 -242
rect 1383 -246 1384 -244
rect 1386 -246 1387 -244
rect 1415 -231 1419 -219
rect 1415 -233 1416 -231
rect 1418 -233 1419 -231
rect 1415 -239 1419 -233
rect 1383 -251 1387 -246
rect 1414 -241 1419 -239
rect 1414 -243 1415 -241
rect 1417 -243 1419 -241
rect 1414 -248 1419 -243
rect 1369 -254 1371 -252
rect 1358 -256 1371 -254
rect 1358 -258 1368 -256
rect 1370 -258 1371 -256
rect 1367 -259 1371 -258
rect 1414 -250 1415 -248
rect 1417 -250 1419 -248
rect 1414 -252 1419 -250
rect 1423 -215 1428 -213
rect 1423 -217 1425 -215
rect 1427 -217 1428 -215
rect 1423 -219 1428 -217
rect 1423 -223 1427 -219
rect 1423 -225 1424 -223
rect 1426 -225 1427 -223
rect 1423 -241 1427 -225
rect 1502 -215 1508 -214
rect 1502 -217 1503 -215
rect 1505 -217 1508 -215
rect 1502 -218 1508 -217
rect 1423 -243 1428 -241
rect 1423 -245 1425 -243
rect 1427 -245 1428 -243
rect 1423 -250 1428 -245
rect 1451 -231 1459 -229
rect 1471 -230 1475 -221
rect 1451 -233 1452 -231
rect 1454 -233 1459 -231
rect 1451 -235 1459 -233
rect 1469 -231 1484 -230
rect 1469 -233 1471 -231
rect 1473 -233 1474 -231
rect 1476 -233 1478 -231
rect 1480 -233 1484 -231
rect 1469 -234 1484 -233
rect 1454 -238 1459 -235
rect 1504 -231 1508 -218
rect 1504 -233 1505 -231
rect 1507 -233 1508 -231
rect 1454 -239 1492 -238
rect 1454 -241 1468 -239
rect 1470 -241 1492 -239
rect 1454 -242 1492 -241
rect 1504 -238 1508 -233
rect 1502 -240 1508 -238
rect 1502 -242 1503 -240
rect 1505 -242 1508 -240
rect 1502 -247 1508 -242
rect 1502 -249 1503 -247
rect 1505 -249 1508 -247
rect 1423 -252 1425 -250
rect 1427 -252 1428 -250
rect 1423 -254 1428 -252
rect 1502 -251 1508 -249
rect 1512 -215 1518 -214
rect 1512 -217 1515 -215
rect 1517 -217 1518 -215
rect 1512 -218 1518 -217
rect 1592 -214 1599 -213
rect 1592 -215 1596 -214
rect 1592 -217 1593 -215
rect 1595 -216 1596 -215
rect 1598 -216 1599 -214
rect 1595 -217 1599 -216
rect 1512 -238 1516 -218
rect 1545 -223 1549 -221
rect 1545 -225 1546 -223
rect 1548 -225 1549 -223
rect 1512 -240 1518 -238
rect 1512 -242 1515 -240
rect 1517 -242 1518 -240
rect 1512 -244 1518 -242
rect 1512 -246 1515 -244
rect 1517 -246 1518 -244
rect 1512 -247 1518 -246
rect 1512 -249 1515 -247
rect 1517 -249 1518 -247
rect 1512 -251 1518 -249
rect 1545 -230 1549 -225
rect 1592 -219 1599 -217
rect 1536 -231 1551 -230
rect 1536 -233 1540 -231
rect 1542 -233 1547 -231
rect 1549 -233 1551 -231
rect 1536 -234 1551 -233
rect 1561 -231 1569 -229
rect 1561 -233 1566 -231
rect 1568 -233 1569 -231
rect 1561 -235 1569 -233
rect 1561 -236 1566 -235
rect 1561 -238 1563 -236
rect 1565 -238 1566 -236
rect 1528 -242 1566 -238
rect 1593 -241 1597 -219
rect 1602 -225 1606 -224
rect 1602 -227 1603 -225
rect 1605 -227 1606 -225
rect 1602 -230 1606 -227
rect 1602 -231 1623 -230
rect 1602 -233 1617 -231
rect 1619 -233 1623 -231
rect 1602 -234 1623 -233
rect 1633 -222 1638 -220
rect 1633 -224 1634 -222
rect 1636 -224 1638 -222
rect 1633 -226 1638 -224
rect 1592 -243 1597 -241
rect 1592 -245 1593 -243
rect 1595 -245 1597 -243
rect 1592 -250 1597 -245
rect 1592 -252 1593 -250
rect 1595 -252 1597 -250
rect 1602 -240 1607 -238
rect 1609 -240 1623 -238
rect 1602 -242 1623 -240
rect 1602 -244 1606 -242
rect 1602 -246 1603 -244
rect 1605 -246 1606 -244
rect 1602 -251 1606 -246
rect 1592 -254 1597 -252
rect 1634 -245 1638 -226
rect 1657 -230 1662 -221
rect 1674 -217 1686 -213
rect 1674 -219 1682 -217
rect 1684 -219 1686 -217
rect 1657 -231 1671 -230
rect 1657 -233 1665 -231
rect 1667 -233 1671 -231
rect 1657 -234 1671 -233
rect 1636 -247 1638 -245
rect 1634 -252 1638 -247
rect 1650 -239 1663 -238
rect 1650 -241 1655 -239
rect 1657 -241 1663 -239
rect 1650 -242 1663 -241
rect 1650 -244 1654 -242
rect 1650 -246 1651 -244
rect 1653 -246 1654 -244
rect 1682 -231 1686 -219
rect 1682 -233 1683 -231
rect 1685 -233 1686 -231
rect 1682 -239 1686 -233
rect 1650 -251 1654 -246
rect 1681 -241 1686 -239
rect 1681 -243 1682 -241
rect 1684 -243 1686 -241
rect 1681 -248 1686 -243
rect 1636 -254 1638 -252
rect 1625 -256 1638 -254
rect 1625 -258 1635 -256
rect 1637 -258 1638 -256
rect 1634 -259 1638 -258
rect 1681 -250 1682 -248
rect 1684 -250 1686 -248
rect 1681 -252 1686 -250
rect 1690 -215 1695 -213
rect 1690 -217 1692 -215
rect 1694 -217 1695 -215
rect 1690 -219 1695 -217
rect 1690 -223 1694 -219
rect 1690 -225 1691 -223
rect 1693 -225 1694 -223
rect 1690 -241 1694 -225
rect 1769 -215 1775 -214
rect 1769 -217 1770 -215
rect 1772 -217 1775 -215
rect 1769 -218 1775 -217
rect 1690 -243 1695 -241
rect 1690 -245 1692 -243
rect 1694 -245 1695 -243
rect 1690 -250 1695 -245
rect 1718 -231 1726 -229
rect 1738 -230 1742 -221
rect 1718 -233 1719 -231
rect 1721 -233 1726 -231
rect 1718 -235 1726 -233
rect 1736 -231 1751 -230
rect 1736 -233 1738 -231
rect 1740 -233 1741 -231
rect 1743 -233 1745 -231
rect 1747 -233 1751 -231
rect 1736 -234 1751 -233
rect 1721 -238 1726 -235
rect 1771 -231 1775 -218
rect 1771 -233 1772 -231
rect 1774 -233 1775 -231
rect 1721 -239 1759 -238
rect 1721 -241 1735 -239
rect 1737 -241 1759 -239
rect 1721 -242 1759 -241
rect 1771 -238 1775 -233
rect 1769 -240 1775 -238
rect 1769 -242 1770 -240
rect 1772 -242 1775 -240
rect 1769 -247 1775 -242
rect 1769 -249 1770 -247
rect 1772 -249 1775 -247
rect 1690 -252 1692 -250
rect 1694 -252 1695 -250
rect 1690 -254 1695 -252
rect 1769 -251 1775 -249
rect 1779 -215 1785 -214
rect 1779 -217 1782 -215
rect 1784 -217 1785 -215
rect 1779 -218 1785 -217
rect 1859 -214 1866 -213
rect 1859 -215 1863 -214
rect 1859 -217 1860 -215
rect 1862 -216 1863 -215
rect 1865 -216 1866 -214
rect 1862 -217 1866 -216
rect 1948 -215 1972 -214
rect 1779 -238 1783 -218
rect 1812 -223 1816 -221
rect 1812 -225 1813 -223
rect 1815 -225 1816 -223
rect 1779 -240 1785 -238
rect 1779 -242 1782 -240
rect 1784 -242 1785 -240
rect 1779 -244 1785 -242
rect 1779 -246 1782 -244
rect 1784 -246 1785 -244
rect 1779 -247 1785 -246
rect 1779 -249 1782 -247
rect 1784 -249 1785 -247
rect 1779 -251 1785 -249
rect 1812 -230 1816 -225
rect 1859 -219 1866 -217
rect 1948 -217 1950 -215
rect 1952 -217 1972 -215
rect 1948 -218 1972 -217
rect 1803 -231 1818 -230
rect 1803 -233 1807 -231
rect 1809 -233 1814 -231
rect 1816 -233 1818 -231
rect 1803 -234 1818 -233
rect 1828 -231 1836 -229
rect 1828 -233 1833 -231
rect 1835 -233 1836 -231
rect 1828 -235 1836 -233
rect 1828 -236 1833 -235
rect 1828 -238 1830 -236
rect 1832 -238 1833 -236
rect 1795 -242 1833 -238
rect 1860 -241 1864 -219
rect 1869 -225 1873 -224
rect 1869 -227 1870 -225
rect 1872 -227 1873 -225
rect 1869 -230 1873 -227
rect 1869 -231 1890 -230
rect 1869 -233 1884 -231
rect 1886 -233 1890 -231
rect 1869 -234 1890 -233
rect 1900 -222 1905 -220
rect 1900 -224 1901 -222
rect 1903 -224 1905 -222
rect 1900 -226 1905 -224
rect 1859 -243 1864 -241
rect 1859 -245 1860 -243
rect 1862 -245 1864 -243
rect 1859 -250 1864 -245
rect 1859 -252 1860 -250
rect 1862 -252 1864 -250
rect 1869 -240 1874 -238
rect 1876 -240 1890 -238
rect 1869 -242 1890 -240
rect 1869 -244 1873 -242
rect 1869 -246 1870 -244
rect 1872 -246 1873 -244
rect 1869 -251 1873 -246
rect 1859 -254 1864 -252
rect 1901 -245 1905 -226
rect 1920 -222 1933 -221
rect 1920 -224 1925 -222
rect 1927 -224 1933 -222
rect 1920 -226 1933 -224
rect 1920 -227 1930 -226
rect 1928 -228 1930 -227
rect 1932 -228 1933 -226
rect 1903 -247 1905 -245
rect 1901 -252 1905 -247
rect 1903 -254 1905 -252
rect 1892 -256 1905 -254
rect 1892 -258 1902 -256
rect 1904 -258 1905 -256
rect 1901 -259 1905 -258
rect 1912 -239 1917 -237
rect 1912 -241 1914 -239
rect 1916 -241 1917 -239
rect 1912 -253 1917 -241
rect 1928 -235 1933 -228
rect 1912 -259 1924 -253
rect 1968 -239 1972 -218
rect 1968 -241 1969 -239
rect 1971 -241 1972 -239
rect 1968 -246 1972 -241
rect 1956 -248 1972 -246
rect 1956 -250 1958 -248
rect 1960 -250 1972 -248
rect 1956 -251 1972 -250
rect 1976 -215 1981 -213
rect 1976 -217 1978 -215
rect 1980 -217 1981 -215
rect 1976 -219 1981 -217
rect 1976 -223 1980 -219
rect 1976 -225 1977 -223
rect 1979 -225 1980 -223
rect 1976 -241 1980 -225
rect 2055 -215 2061 -214
rect 2055 -217 2056 -215
rect 2058 -217 2061 -215
rect 2055 -218 2061 -217
rect 1976 -243 1981 -241
rect 1976 -245 1978 -243
rect 1980 -245 1981 -243
rect 1976 -250 1981 -245
rect 2004 -231 2012 -229
rect 2024 -230 2028 -221
rect 2004 -233 2005 -231
rect 2007 -233 2012 -231
rect 2004 -235 2012 -233
rect 2022 -231 2037 -230
rect 2022 -233 2024 -231
rect 2026 -233 2031 -231
rect 2033 -233 2037 -231
rect 2022 -234 2037 -233
rect 2007 -238 2012 -235
rect 2057 -231 2061 -218
rect 2057 -233 2058 -231
rect 2060 -233 2061 -231
rect 2007 -239 2045 -238
rect 2007 -241 2018 -239
rect 2020 -241 2045 -239
rect 2007 -242 2045 -241
rect 2057 -238 2061 -233
rect 2055 -240 2061 -238
rect 2055 -242 2056 -240
rect 2058 -242 2061 -240
rect 2055 -247 2061 -242
rect 2055 -249 2056 -247
rect 2058 -249 2061 -247
rect 1976 -252 1978 -250
rect 1980 -252 1981 -250
rect 1976 -254 1981 -252
rect 2055 -251 2061 -249
rect 2065 -215 2071 -214
rect 2065 -217 2068 -215
rect 2070 -217 2071 -215
rect 2065 -218 2071 -217
rect 2145 -214 2152 -213
rect 2145 -215 2149 -214
rect 2145 -217 2146 -215
rect 2148 -216 2149 -215
rect 2151 -216 2152 -214
rect 2148 -217 2152 -216
rect 2065 -238 2069 -218
rect 2098 -223 2102 -221
rect 2098 -225 2099 -223
rect 2101 -225 2102 -223
rect 2065 -240 2071 -238
rect 2065 -242 2068 -240
rect 2070 -242 2071 -240
rect 2065 -244 2071 -242
rect 2065 -246 2068 -244
rect 2070 -246 2071 -244
rect 2065 -247 2071 -246
rect 2065 -249 2068 -247
rect 2070 -249 2071 -247
rect 2065 -251 2071 -249
rect 2098 -230 2102 -225
rect 2145 -219 2150 -217
rect 2089 -231 2104 -230
rect 2089 -233 2093 -231
rect 2095 -233 2100 -231
rect 2102 -233 2104 -231
rect 2089 -234 2104 -233
rect 2114 -231 2122 -229
rect 2114 -233 2119 -231
rect 2121 -233 2122 -231
rect 2114 -235 2122 -233
rect 2114 -236 2119 -235
rect 2114 -238 2116 -236
rect 2118 -238 2119 -236
rect 2081 -242 2119 -238
rect 2146 -241 2150 -219
rect 2155 -225 2159 -221
rect 2155 -227 2156 -225
rect 2158 -227 2159 -225
rect 2155 -230 2159 -227
rect 2155 -231 2176 -230
rect 2155 -233 2170 -231
rect 2172 -233 2176 -231
rect 2155 -234 2176 -233
rect 2186 -222 2191 -220
rect 2186 -224 2187 -222
rect 2189 -224 2191 -222
rect 2186 -226 2191 -224
rect 2145 -243 2150 -241
rect 2145 -245 2146 -243
rect 2148 -245 2150 -243
rect 2145 -250 2150 -245
rect 2145 -252 2146 -250
rect 2148 -252 2150 -250
rect 2155 -240 2160 -238
rect 2162 -240 2176 -238
rect 2155 -242 2176 -240
rect 2155 -244 2159 -242
rect 2155 -246 2156 -244
rect 2158 -246 2159 -244
rect 2187 -228 2191 -226
rect 2187 -230 2188 -228
rect 2190 -230 2191 -228
rect 2155 -251 2159 -246
rect 2145 -254 2150 -252
rect 2187 -245 2191 -230
rect 2255 -215 2259 -213
rect 2254 -217 2259 -215
rect 2254 -219 2255 -217
rect 2257 -219 2259 -217
rect 2254 -221 2259 -219
rect 2206 -223 2219 -222
rect 2206 -225 2210 -223
rect 2212 -225 2219 -223
rect 2206 -226 2219 -225
rect 2213 -231 2219 -226
rect 2213 -233 2214 -231
rect 2216 -233 2219 -231
rect 2213 -235 2219 -233
rect 2239 -236 2243 -229
rect 2239 -237 2241 -236
rect 2231 -238 2241 -237
rect 2231 -240 2243 -238
rect 2231 -242 2236 -240
rect 2238 -242 2243 -240
rect 2231 -243 2243 -242
rect 2189 -247 2191 -245
rect 2187 -252 2191 -247
rect 2189 -254 2191 -252
rect 2178 -258 2191 -254
rect 2187 -259 2191 -258
rect 2199 -250 2212 -246
rect 2199 -251 2204 -250
rect 2199 -253 2201 -251
rect 2203 -253 2204 -251
rect 2199 -259 2204 -253
rect 2255 -254 2259 -221
rect 2323 -215 2327 -213
rect 2322 -217 2327 -215
rect 2322 -219 2323 -217
rect 2325 -219 2327 -217
rect 2322 -221 2327 -219
rect 2274 -223 2287 -222
rect 2274 -225 2276 -223
rect 2278 -225 2287 -223
rect 2274 -226 2287 -225
rect 2281 -231 2287 -226
rect 2281 -233 2282 -231
rect 2284 -233 2287 -231
rect 2281 -235 2287 -233
rect 2307 -236 2311 -229
rect 2307 -237 2309 -236
rect 2299 -238 2309 -237
rect 2299 -240 2300 -238
rect 2302 -240 2311 -238
rect 2299 -243 2311 -240
rect 2246 -255 2259 -254
rect 2246 -257 2255 -255
rect 2257 -257 2259 -255
rect 2246 -258 2259 -257
rect 2267 -250 2280 -246
rect 2267 -251 2272 -250
rect 2267 -253 2269 -251
rect 2271 -253 2272 -251
rect 2267 -259 2272 -253
rect 2323 -254 2327 -221
rect 2314 -255 2327 -254
rect 2314 -257 2323 -255
rect 2325 -257 2327 -255
rect 2314 -258 2327 -257
rect 4 -265 2331 -264
rect 4 -267 39 -265
rect 41 -267 79 -265
rect 81 -267 298 -265
rect 300 -267 346 -265
rect 348 -267 565 -265
rect 567 -267 613 -265
rect 615 -267 832 -265
rect 834 -267 880 -265
rect 882 -267 1099 -265
rect 1101 -267 1147 -265
rect 1149 -267 1366 -265
rect 1368 -267 1414 -265
rect 1416 -267 1633 -265
rect 1635 -267 1681 -265
rect 1683 -267 1900 -265
rect 1902 -267 1948 -265
rect 1950 -267 2186 -265
rect 2188 -267 2328 -265
rect 2330 -267 2331 -265
rect 4 -272 2331 -267
<< alu2 >>
rect 2319 303 2327 304
rect 2319 301 2320 303
rect 2322 301 2324 303
rect 2326 301 2327 303
rect 2319 300 2327 301
rect 1928 290 2095 291
rect 1928 288 1929 290
rect 1931 288 2092 290
rect 2094 288 2095 290
rect 1928 287 2095 288
rect 183 282 271 283
rect 183 280 268 282
rect 270 280 271 282
rect 183 279 271 280
rect 450 282 538 283
rect 450 280 535 282
rect 537 280 538 282
rect 450 279 538 280
rect 717 282 805 283
rect 717 280 802 282
rect 804 280 805 282
rect 717 279 805 280
rect 984 282 1072 283
rect 984 280 1069 282
rect 1071 280 1072 282
rect 984 279 1072 280
rect 1251 282 1339 283
rect 1251 280 1336 282
rect 1338 280 1339 282
rect 1251 279 1339 280
rect 1518 282 1606 283
rect 1518 280 1603 282
rect 1605 280 1606 282
rect 1518 279 1606 280
rect 1785 282 1873 283
rect 1785 280 1870 282
rect 1872 280 1873 282
rect 1785 279 1873 280
rect 2075 279 2151 283
rect 179 278 187 279
rect 2 276 12 277
rect 2 274 3 276
rect 5 274 9 276
rect 11 274 12 276
rect 179 276 180 278
rect 182 276 187 278
rect 179 275 187 276
rect 446 278 454 279
rect 446 276 447 278
rect 449 276 454 278
rect 446 275 454 276
rect 713 278 721 279
rect 713 276 714 278
rect 716 276 721 278
rect 713 275 721 276
rect 980 278 988 279
rect 980 276 981 278
rect 983 276 988 278
rect 980 275 988 276
rect 1247 278 1255 279
rect 1247 276 1248 278
rect 1250 276 1255 278
rect 1247 275 1255 276
rect 1514 278 1522 279
rect 1514 276 1515 278
rect 1517 276 1522 278
rect 1514 275 1522 276
rect 1781 278 1789 279
rect 1781 276 1782 278
rect 1784 276 1789 278
rect 1781 275 1789 276
rect 2067 278 2079 279
rect 2067 276 2068 278
rect 2070 276 2079 278
rect 2067 275 2079 276
rect 2147 278 2159 279
rect 2147 276 2156 278
rect 2158 276 2159 278
rect 2147 275 2159 276
rect 262 274 266 275
rect 2299 274 2307 275
rect 2 273 12 274
rect 45 273 124 274
rect 45 271 121 273
rect 123 271 124 273
rect 40 270 124 271
rect 209 273 217 274
rect 209 271 210 273
rect 212 271 213 273
rect 215 271 217 273
rect 209 270 217 271
rect 258 273 263 274
rect 258 271 259 273
rect 261 272 263 273
rect 265 272 266 274
rect 261 271 266 272
rect 258 270 266 271
rect 351 273 391 274
rect 351 271 352 273
rect 354 271 388 273
rect 390 271 391 273
rect 351 270 391 271
rect 476 273 484 274
rect 476 271 477 273
rect 479 271 480 273
rect 482 271 484 273
rect 476 270 484 271
rect 525 273 533 274
rect 525 271 526 273
rect 528 271 530 273
rect 532 271 533 273
rect 525 270 533 271
rect 618 273 658 274
rect 618 271 619 273
rect 621 271 655 273
rect 657 271 658 273
rect 618 270 658 271
rect 743 273 751 274
rect 743 271 744 273
rect 746 271 747 273
rect 749 271 751 273
rect 743 270 751 271
rect 885 273 925 274
rect 885 271 886 273
rect 888 271 922 273
rect 924 271 925 273
rect 885 270 925 271
rect 1010 273 1018 274
rect 1010 271 1011 273
rect 1013 271 1014 273
rect 1016 271 1018 273
rect 1010 270 1018 271
rect 1152 273 1192 274
rect 1152 271 1153 273
rect 1155 271 1189 273
rect 1191 271 1192 273
rect 1152 270 1192 271
rect 1277 273 1285 274
rect 1277 271 1278 273
rect 1280 271 1281 273
rect 1283 271 1285 273
rect 1277 270 1285 271
rect 1419 273 1459 274
rect 1419 271 1420 273
rect 1422 271 1456 273
rect 1458 271 1459 273
rect 1419 270 1459 271
rect 1544 273 1552 274
rect 1544 271 1545 273
rect 1547 271 1548 273
rect 1550 271 1552 273
rect 1544 270 1552 271
rect 1686 273 1726 274
rect 1686 271 1687 273
rect 1689 271 1723 273
rect 1725 271 1726 273
rect 1686 270 1726 271
rect 1811 273 1819 274
rect 1811 271 1812 273
rect 1814 271 1815 273
rect 1817 271 1819 273
rect 1811 270 1819 271
rect 1860 273 1864 274
rect 1860 271 1861 273
rect 1863 271 1864 273
rect 1860 270 1864 271
rect 1968 273 2021 274
rect 1968 271 1969 273
rect 1971 271 2018 273
rect 2020 271 2021 273
rect 1968 270 2021 271
rect 2091 273 2103 274
rect 2091 271 2092 273
rect 2094 271 2100 273
rect 2102 271 2103 273
rect 2091 270 2103 271
rect 2192 273 2239 274
rect 2192 271 2193 273
rect 2195 271 2236 273
rect 2238 271 2239 273
rect 2299 272 2300 274
rect 2302 272 2304 274
rect 2306 272 2307 274
rect 2299 271 2307 272
rect 2192 270 2239 271
rect 40 268 41 270
rect 43 268 49 270
rect 40 267 49 268
rect 80 265 142 266
rect 80 263 81 265
rect 83 263 139 265
rect 141 263 142 265
rect 80 262 142 263
rect 169 265 272 266
rect 169 263 170 265
rect 172 263 268 265
rect 270 263 272 265
rect 169 262 272 263
rect 347 265 409 266
rect 347 263 348 265
rect 350 263 406 265
rect 408 263 409 265
rect 347 262 409 263
rect 436 265 539 266
rect 436 263 437 265
rect 439 263 535 265
rect 537 263 539 265
rect 436 262 539 263
rect 614 265 676 266
rect 614 263 615 265
rect 617 263 673 265
rect 675 263 676 265
rect 614 262 676 263
rect 703 265 806 266
rect 703 263 704 265
rect 706 263 802 265
rect 804 263 806 265
rect 703 262 806 263
rect 881 265 943 266
rect 881 263 882 265
rect 884 263 940 265
rect 942 263 943 265
rect 881 262 943 263
rect 970 265 1073 266
rect 970 263 971 265
rect 973 263 1069 265
rect 1071 263 1073 265
rect 970 262 1073 263
rect 1148 265 1210 266
rect 1148 263 1149 265
rect 1151 263 1207 265
rect 1209 263 1210 265
rect 1148 262 1210 263
rect 1237 265 1340 266
rect 1237 263 1238 265
rect 1240 263 1336 265
rect 1338 263 1340 265
rect 1237 262 1340 263
rect 1415 265 1477 266
rect 1415 263 1416 265
rect 1418 263 1474 265
rect 1476 263 1477 265
rect 1415 262 1477 263
rect 1504 265 1607 266
rect 1504 263 1505 265
rect 1507 263 1603 265
rect 1605 263 1607 265
rect 1504 262 1607 263
rect 1682 265 1744 266
rect 1682 263 1683 265
rect 1685 263 1741 265
rect 1743 263 1744 265
rect 1682 262 1744 263
rect 1771 265 1874 266
rect 1771 263 1772 265
rect 1774 263 1870 265
rect 1872 263 1874 265
rect 1771 262 1874 263
rect 2057 265 2160 266
rect 2057 263 2058 265
rect 2060 263 2156 265
rect 2158 263 2160 265
rect 2057 262 2160 263
rect 299 261 307 262
rect 44 259 60 260
rect 44 257 45 259
rect 47 257 57 259
rect 59 257 60 259
rect 299 259 300 261
rect 302 259 304 261
rect 306 259 307 261
rect 566 261 574 262
rect 299 258 307 259
rect 311 259 327 260
rect 44 255 60 257
rect 88 257 214 258
rect 88 255 89 257
rect 91 255 211 257
rect 213 255 214 257
rect 311 257 312 259
rect 314 257 324 259
rect 326 257 327 259
rect 566 259 567 261
rect 569 259 571 261
rect 573 259 574 261
rect 833 261 841 262
rect 566 258 574 259
rect 578 259 594 260
rect 311 255 327 257
rect 355 257 481 258
rect 355 255 356 257
rect 358 255 478 257
rect 480 255 481 257
rect 578 257 579 259
rect 581 257 591 259
rect 593 257 594 259
rect 833 259 834 261
rect 836 259 838 261
rect 840 259 841 261
rect 1100 261 1108 262
rect 833 258 841 259
rect 845 259 861 260
rect 578 255 594 257
rect 622 257 748 258
rect 622 255 623 257
rect 625 255 745 257
rect 747 255 748 257
rect 88 254 214 255
rect 355 254 481 255
rect 622 254 748 255
rect 792 257 800 258
rect 792 255 793 257
rect 795 255 797 257
rect 799 255 800 257
rect 845 257 846 259
rect 848 257 858 259
rect 860 257 861 259
rect 1100 259 1101 261
rect 1103 259 1105 261
rect 1107 259 1108 261
rect 1367 261 1375 262
rect 1100 258 1108 259
rect 1112 259 1128 260
rect 845 255 861 257
rect 889 257 1015 258
rect 889 255 890 257
rect 892 255 1012 257
rect 1014 255 1015 257
rect 792 254 800 255
rect 889 254 1015 255
rect 1059 257 1067 258
rect 1059 255 1060 257
rect 1062 255 1064 257
rect 1066 255 1067 257
rect 1112 257 1113 259
rect 1115 257 1125 259
rect 1127 257 1128 259
rect 1367 259 1368 261
rect 1370 259 1372 261
rect 1374 259 1375 261
rect 1634 261 1642 262
rect 1367 258 1375 259
rect 1379 259 1395 260
rect 1112 255 1128 257
rect 1156 257 1282 258
rect 1156 255 1157 257
rect 1159 255 1279 257
rect 1281 255 1282 257
rect 1379 257 1380 259
rect 1382 257 1392 259
rect 1394 257 1395 259
rect 1634 259 1635 261
rect 1637 259 1639 261
rect 1641 259 1642 261
rect 1901 261 1909 262
rect 1634 258 1642 259
rect 1646 259 1662 260
rect 1379 255 1395 257
rect 1423 257 1549 258
rect 1423 255 1424 257
rect 1426 255 1546 257
rect 1548 255 1549 257
rect 1646 257 1647 259
rect 1649 257 1659 259
rect 1661 257 1662 259
rect 1901 259 1902 261
rect 1904 259 1906 261
rect 1908 259 1909 261
rect 1901 258 1909 259
rect 2187 261 2195 262
rect 2187 259 2188 261
rect 2190 259 2192 261
rect 2194 259 2195 261
rect 2187 258 2195 259
rect 1646 255 1662 257
rect 1690 257 1816 258
rect 1976 257 2102 258
rect 1690 255 1691 257
rect 1693 255 1813 257
rect 1815 255 1816 257
rect 1059 254 1067 255
rect 1156 254 1282 255
rect 1326 254 1330 255
rect 1423 254 1549 255
rect 1593 254 1601 255
rect 1690 254 1816 255
rect 1924 256 1932 257
rect 1924 254 1925 256
rect 1927 254 1929 256
rect 1931 254 1932 256
rect 1976 255 1977 257
rect 1979 255 2099 257
rect 2101 255 2102 257
rect 1976 254 2102 255
rect 2146 257 2150 258
rect 2146 255 2147 257
rect 2149 255 2150 257
rect 2146 254 2150 255
rect 2207 257 2211 258
rect 2207 255 2208 257
rect 2210 255 2211 257
rect 2207 254 2211 255
rect 1326 252 1327 254
rect 1329 252 1330 254
rect 1326 249 1330 252
rect 1593 252 1594 254
rect 1596 252 1601 254
rect 1924 253 1932 254
rect 1593 251 1601 252
rect 1597 250 1601 251
rect 2146 250 2211 254
rect 2263 257 2279 258
rect 2263 255 2276 257
rect 2278 255 2279 257
rect 2263 254 2279 255
rect 1326 248 1334 249
rect 1326 246 1331 248
rect 1333 246 1334 248
rect 1597 248 1598 250
rect 1600 248 1601 250
rect 1597 247 1601 248
rect 1326 245 1334 246
rect 212 236 219 237
rect 212 234 213 236
rect 215 234 216 236
rect 218 234 219 236
rect 212 233 219 234
rect 479 236 486 237
rect 479 234 480 236
rect 482 234 483 236
rect 485 234 486 236
rect 479 233 486 234
rect 746 236 753 237
rect 746 234 747 236
rect 749 234 750 236
rect 752 234 753 236
rect 746 233 753 234
rect 1013 236 1020 237
rect 1013 234 1014 236
rect 1016 234 1017 236
rect 1019 234 1020 236
rect 1013 233 1020 234
rect 1280 236 1287 237
rect 1280 234 1281 236
rect 1283 234 1284 236
rect 1286 234 1287 236
rect 1280 233 1287 234
rect 1547 236 1554 237
rect 1547 234 1548 236
rect 1550 234 1551 236
rect 1553 234 1554 236
rect 1547 233 1554 234
rect 1814 236 1821 237
rect 1814 234 1815 236
rect 1817 234 1818 236
rect 1820 234 1821 236
rect 1814 233 1821 234
rect 2263 226 2267 254
rect 2263 224 2264 226
rect 2266 224 2267 226
rect 2263 223 2267 224
rect 2275 233 2279 234
rect 2275 231 2276 233
rect 2278 231 2279 233
rect 260 218 355 219
rect 260 216 261 218
rect 263 216 352 218
rect 354 216 355 218
rect 260 215 355 216
rect 527 218 622 219
rect 527 216 528 218
rect 530 216 619 218
rect 621 216 622 218
rect 527 215 622 216
rect 794 218 889 219
rect 794 216 795 218
rect 797 216 886 218
rect 888 216 889 218
rect 794 215 889 216
rect 1061 218 1156 219
rect 1061 216 1062 218
rect 1064 216 1153 218
rect 1155 216 1156 218
rect 1061 215 1156 216
rect 1328 218 1423 219
rect 1328 216 1329 218
rect 1331 216 1420 218
rect 1422 216 1423 218
rect 1328 215 1423 216
rect 1595 218 1690 219
rect 1595 216 1596 218
rect 1598 216 1687 218
rect 1689 216 1690 218
rect 1595 215 1690 216
rect 1862 218 1884 219
rect 1862 216 1863 218
rect 1865 216 1881 218
rect 1883 216 1884 218
rect 1862 215 1884 216
rect 2148 218 2167 219
rect 2148 216 2149 218
rect 2151 216 2167 218
rect 2148 215 2167 216
rect 1924 210 1932 211
rect 2163 210 2167 215
rect 88 209 214 210
rect 88 207 89 209
rect 91 207 211 209
rect 213 207 214 209
rect 355 209 481 210
rect 88 206 214 207
rect 218 207 271 208
rect 2 205 20 206
rect 2 203 3 205
rect 5 203 17 205
rect 19 203 20 205
rect 2 202 20 203
rect 218 205 268 207
rect 270 205 271 207
rect 355 207 356 209
rect 358 207 478 209
rect 480 207 481 209
rect 622 209 748 210
rect 355 206 481 207
rect 485 207 538 208
rect 218 204 271 205
rect 485 205 535 207
rect 537 205 538 207
rect 622 207 623 209
rect 625 207 745 209
rect 747 207 748 209
rect 889 209 1015 210
rect 622 206 748 207
rect 752 207 805 208
rect 485 204 538 205
rect 752 205 802 207
rect 804 205 805 207
rect 889 207 890 209
rect 892 207 1012 209
rect 1014 207 1015 209
rect 1156 209 1282 210
rect 889 206 1015 207
rect 1019 207 1072 208
rect 752 204 805 205
rect 1019 205 1069 207
rect 1071 205 1072 207
rect 1156 207 1157 209
rect 1159 207 1279 209
rect 1281 207 1282 209
rect 1423 209 1549 210
rect 1156 206 1282 207
rect 1286 207 1339 208
rect 1019 204 1072 205
rect 1286 205 1336 207
rect 1338 205 1339 207
rect 1423 207 1424 209
rect 1426 207 1546 209
rect 1548 207 1549 209
rect 1690 209 1816 210
rect 1423 206 1549 207
rect 1553 207 1606 208
rect 1286 204 1339 205
rect 1553 205 1603 207
rect 1605 205 1606 207
rect 1690 207 1691 209
rect 1693 207 1813 209
rect 1815 207 1816 209
rect 1924 208 1925 210
rect 1927 208 1929 210
rect 1931 208 1932 210
rect 1690 206 1816 207
rect 1820 207 1873 208
rect 1924 207 1932 208
rect 1976 209 2102 210
rect 1976 207 1977 209
rect 1979 207 2099 209
rect 2101 207 2102 209
rect 2163 209 2213 210
rect 1553 204 1606 205
rect 1820 205 1870 207
rect 1872 205 1873 207
rect 1976 206 2102 207
rect 2106 207 2159 208
rect 1820 204 1873 205
rect 2106 205 2156 207
rect 2158 205 2159 207
rect 2163 207 2210 209
rect 2212 207 2213 209
rect 2163 206 2213 207
rect 2275 209 2279 231
rect 2310 229 2318 230
rect 2310 227 2311 229
rect 2313 227 2315 229
rect 2317 227 2318 229
rect 2310 226 2318 227
rect 2275 207 2276 209
rect 2278 207 2279 209
rect 2275 206 2279 207
rect 2106 204 2159 205
rect 218 202 222 204
rect 485 202 489 204
rect 752 202 756 204
rect 1019 202 1023 204
rect 1286 202 1290 204
rect 1553 202 1557 204
rect 1820 202 1824 204
rect 2106 202 2110 204
rect 80 201 142 202
rect 80 199 81 201
rect 83 199 139 201
rect 141 199 142 201
rect 80 198 142 199
rect 169 201 222 202
rect 169 199 170 201
rect 172 199 222 201
rect 169 198 222 199
rect 347 201 409 202
rect 347 199 348 201
rect 350 199 406 201
rect 408 199 409 201
rect 347 198 409 199
rect 436 201 489 202
rect 436 199 437 201
rect 439 199 489 201
rect 436 198 489 199
rect 614 201 676 202
rect 614 199 615 201
rect 617 199 673 201
rect 675 199 676 201
rect 614 198 676 199
rect 703 201 756 202
rect 703 199 704 201
rect 706 199 756 201
rect 703 198 756 199
rect 881 201 943 202
rect 881 199 882 201
rect 884 199 940 201
rect 942 199 943 201
rect 881 198 943 199
rect 970 201 1023 202
rect 970 199 971 201
rect 973 199 1023 201
rect 970 198 1023 199
rect 1148 201 1210 202
rect 1148 199 1149 201
rect 1151 199 1207 201
rect 1209 199 1210 201
rect 1148 198 1210 199
rect 1237 201 1290 202
rect 1237 199 1238 201
rect 1240 199 1290 201
rect 1237 198 1290 199
rect 1415 201 1477 202
rect 1415 199 1416 201
rect 1418 199 1474 201
rect 1476 199 1477 201
rect 1415 198 1477 199
rect 1504 201 1557 202
rect 1504 199 1505 201
rect 1507 199 1557 201
rect 1504 198 1557 199
rect 1682 201 1744 202
rect 1682 199 1683 201
rect 1685 199 1741 201
rect 1743 199 1744 201
rect 1682 198 1744 199
rect 1771 201 1824 202
rect 1771 199 1772 201
rect 1774 199 1824 201
rect 1771 198 1824 199
rect 2057 201 2110 202
rect 2057 199 2058 201
rect 2060 199 2110 201
rect 2057 198 2110 199
rect 2235 200 2239 201
rect 2235 198 2236 200
rect 2238 198 2239 200
rect 227 196 307 197
rect 227 194 228 196
rect 230 194 304 196
rect 306 194 307 196
rect 494 196 574 197
rect 494 194 495 196
rect 497 194 571 196
rect 573 194 574 196
rect 761 196 841 197
rect 761 194 762 196
rect 764 194 838 196
rect 840 194 841 196
rect 1028 196 1108 197
rect 1028 194 1029 196
rect 1031 194 1105 196
rect 1107 194 1108 196
rect 1295 196 1375 197
rect 1295 194 1296 196
rect 1298 194 1372 196
rect 1374 194 1375 196
rect 1562 196 1642 197
rect 1562 194 1563 196
rect 1565 194 1639 196
rect 1641 194 1642 196
rect 1829 196 1909 197
rect 1829 194 1830 196
rect 1832 194 1906 196
rect 1908 194 1909 196
rect 2115 196 2195 197
rect 2115 194 2116 196
rect 2118 194 2192 196
rect 2194 194 2195 196
rect 40 193 137 194
rect 227 193 307 194
rect 335 193 404 194
rect 494 193 574 194
rect 602 193 671 194
rect 761 193 841 194
rect 869 193 938 194
rect 1028 193 1108 194
rect 1136 193 1205 194
rect 1295 193 1375 194
rect 1403 193 1472 194
rect 1562 193 1642 194
rect 1670 193 1739 194
rect 1829 193 1909 194
rect 1968 193 2021 194
rect 2115 193 2195 194
rect 2235 193 2239 198
rect 40 191 41 193
rect 43 191 134 193
rect 136 191 137 193
rect 40 190 137 191
rect 335 191 336 193
rect 338 191 401 193
rect 403 191 404 193
rect 335 190 404 191
rect 602 191 603 193
rect 605 191 668 193
rect 670 191 671 193
rect 602 190 671 191
rect 869 191 870 193
rect 872 191 935 193
rect 937 191 938 193
rect 869 190 938 191
rect 1136 191 1137 193
rect 1139 191 1202 193
rect 1204 191 1205 193
rect 1136 190 1205 191
rect 1403 191 1404 193
rect 1406 191 1469 193
rect 1471 191 1472 193
rect 1403 190 1472 191
rect 1670 191 1671 193
rect 1673 191 1736 193
rect 1738 191 1739 193
rect 1670 190 1739 191
rect 1968 191 1969 193
rect 1971 191 2018 193
rect 2020 191 2021 193
rect 1968 190 2021 191
rect 2235 191 2236 193
rect 2238 191 2239 193
rect 2299 194 2307 195
rect 2299 192 2300 194
rect 2302 192 2304 194
rect 2306 192 2307 194
rect 2299 191 2307 192
rect 2235 190 2239 191
rect 179 188 271 189
rect 179 186 180 188
rect 182 186 268 188
rect 270 186 271 188
rect 446 188 538 189
rect 446 186 447 188
rect 449 186 535 188
rect 537 186 538 188
rect 713 188 805 189
rect 713 186 714 188
rect 716 186 802 188
rect 804 186 805 188
rect 980 188 1072 189
rect 980 186 981 188
rect 983 186 1069 188
rect 1071 186 1072 188
rect 1247 188 1339 189
rect 1247 186 1248 188
rect 1250 186 1336 188
rect 1338 186 1339 188
rect 1514 188 1606 189
rect 1514 186 1515 188
rect 1517 186 1603 188
rect 1605 186 1606 188
rect 1781 188 1873 189
rect 1781 186 1782 188
rect 1784 186 1870 188
rect 1872 186 1873 188
rect 44 185 52 186
rect 179 185 271 186
rect 311 185 319 186
rect 446 185 538 186
rect 578 185 586 186
rect 713 185 805 186
rect 845 185 853 186
rect 980 185 1072 186
rect 1112 185 1120 186
rect 1247 185 1339 186
rect 1379 185 1387 186
rect 1514 185 1606 186
rect 1646 185 1654 186
rect 1781 185 1873 186
rect 2067 188 2159 189
rect 2067 186 2068 188
rect 2070 186 2156 188
rect 2158 186 2159 188
rect 2067 185 2159 186
rect 44 183 45 185
rect 47 183 49 185
rect 51 183 52 185
rect 44 182 52 183
rect 311 183 312 185
rect 314 183 316 185
rect 318 183 319 185
rect 311 182 319 183
rect 578 183 579 185
rect 581 183 583 185
rect 585 183 586 185
rect 578 182 586 183
rect 845 183 846 185
rect 848 183 850 185
rect 852 183 853 185
rect 845 182 853 183
rect 1112 183 1113 185
rect 1115 183 1117 185
rect 1119 183 1120 185
rect 1112 182 1120 183
rect 1379 183 1380 185
rect 1382 183 1384 185
rect 1386 183 1387 185
rect 1379 182 1387 183
rect 1646 183 1647 185
rect 1649 183 1651 185
rect 1653 183 1654 185
rect 1646 182 1654 183
rect 291 177 295 178
rect 291 175 292 177
rect 294 175 295 177
rect 219 138 271 139
rect 219 136 268 138
rect 270 136 271 138
rect 219 135 271 136
rect 179 134 223 135
rect 2 132 12 133
rect 2 130 3 132
rect 5 130 9 132
rect 11 130 12 132
rect 179 132 180 134
rect 182 132 223 134
rect 179 131 223 132
rect 291 130 295 175
rect 558 177 562 178
rect 558 175 559 177
rect 561 175 562 177
rect 486 138 538 139
rect 486 136 535 138
rect 537 136 538 138
rect 486 135 538 136
rect 446 134 490 135
rect 446 132 447 134
rect 449 132 490 134
rect 446 131 490 132
rect 558 130 562 175
rect 825 177 829 178
rect 825 175 826 177
rect 828 175 829 177
rect 753 138 805 139
rect 753 136 802 138
rect 804 136 805 138
rect 753 135 805 136
rect 713 134 757 135
rect 713 132 714 134
rect 716 132 757 134
rect 713 131 757 132
rect 825 130 829 175
rect 1092 177 1096 178
rect 1092 175 1093 177
rect 1095 175 1096 177
rect 1020 138 1072 139
rect 1020 136 1069 138
rect 1071 136 1072 138
rect 1020 135 1072 136
rect 980 134 1024 135
rect 980 132 981 134
rect 983 132 1024 134
rect 980 131 1024 132
rect 1092 130 1096 175
rect 1359 177 1363 178
rect 1359 175 1360 177
rect 1362 175 1363 177
rect 1287 138 1339 139
rect 1287 136 1336 138
rect 1338 136 1339 138
rect 1287 135 1339 136
rect 1247 134 1291 135
rect 1247 132 1248 134
rect 1250 132 1291 134
rect 1247 131 1291 132
rect 1359 130 1363 175
rect 1626 177 1630 178
rect 1626 175 1627 177
rect 1629 175 1630 177
rect 1554 138 1606 139
rect 1554 136 1603 138
rect 1605 136 1606 138
rect 1554 135 1606 136
rect 1514 134 1558 135
rect 1514 132 1515 134
rect 1517 132 1558 134
rect 1514 131 1558 132
rect 1626 130 1630 175
rect 1893 177 1897 178
rect 1893 175 1894 177
rect 1896 175 1897 177
rect 1821 138 1873 139
rect 1821 136 1870 138
rect 1872 136 1873 138
rect 1821 135 1873 136
rect 1781 134 1825 135
rect 1781 132 1782 134
rect 1784 132 1825 134
rect 1781 131 1825 132
rect 1893 130 1897 175
rect 2179 177 2183 178
rect 2179 175 2180 177
rect 2182 175 2183 177
rect 2107 138 2159 139
rect 2107 136 2156 138
rect 2158 136 2159 138
rect 2107 135 2159 136
rect 2067 134 2111 135
rect 2067 132 2068 134
rect 2070 132 2111 134
rect 2067 131 2111 132
rect 2179 130 2183 175
rect 2319 167 2327 168
rect 2319 165 2320 167
rect 2322 165 2324 167
rect 2326 165 2327 167
rect 2319 164 2327 165
rect 2299 130 2307 131
rect 2 129 12 130
rect 39 129 141 130
rect 39 127 41 129
rect 43 127 138 129
rect 140 127 141 129
rect 39 126 141 127
rect 227 129 295 130
rect 227 127 228 129
rect 230 127 295 129
rect 227 126 295 127
rect 351 129 408 130
rect 351 127 352 129
rect 354 127 405 129
rect 407 127 408 129
rect 351 126 408 127
rect 494 129 562 130
rect 494 127 495 129
rect 497 127 562 129
rect 494 126 562 127
rect 618 129 675 130
rect 618 127 619 129
rect 621 127 672 129
rect 674 127 675 129
rect 618 126 675 127
rect 761 129 829 130
rect 761 127 762 129
rect 764 127 829 129
rect 761 126 829 127
rect 885 129 942 130
rect 885 127 886 129
rect 888 127 939 129
rect 941 127 942 129
rect 885 126 942 127
rect 1028 129 1096 130
rect 1028 127 1029 129
rect 1031 127 1096 129
rect 1028 126 1096 127
rect 1152 129 1209 130
rect 1152 127 1153 129
rect 1155 127 1206 129
rect 1208 127 1209 129
rect 1152 126 1209 127
rect 1295 129 1363 130
rect 1295 127 1296 129
rect 1298 127 1363 129
rect 1295 126 1363 127
rect 1419 129 1476 130
rect 1419 127 1420 129
rect 1422 127 1473 129
rect 1475 127 1476 129
rect 1419 126 1476 127
rect 1562 129 1630 130
rect 1562 127 1563 129
rect 1565 127 1630 129
rect 1562 126 1630 127
rect 1686 129 1743 130
rect 1686 127 1687 129
rect 1689 127 1740 129
rect 1742 127 1743 129
rect 1686 126 1743 127
rect 1829 129 1897 130
rect 1829 127 1830 129
rect 1832 127 1897 129
rect 1829 126 1897 127
rect 1968 129 2021 130
rect 1968 127 1969 129
rect 1971 127 2018 129
rect 2020 127 2021 129
rect 1968 126 2021 127
rect 2115 129 2183 130
rect 2115 127 2116 129
rect 2118 127 2183 129
rect 2115 126 2183 127
rect 2227 129 2239 130
rect 2227 127 2228 129
rect 2230 127 2236 129
rect 2238 127 2239 129
rect 2299 128 2300 130
rect 2302 128 2304 130
rect 2306 128 2307 130
rect 2299 127 2307 128
rect 2227 126 2239 127
rect 80 121 143 122
rect 80 119 81 121
rect 83 119 140 121
rect 142 119 143 121
rect 80 118 143 119
rect 169 121 272 122
rect 169 119 170 121
rect 172 119 268 121
rect 270 119 272 121
rect 169 118 272 119
rect 347 121 410 122
rect 347 119 348 121
rect 350 119 407 121
rect 409 119 410 121
rect 347 118 410 119
rect 436 121 539 122
rect 436 119 437 121
rect 439 119 535 121
rect 537 119 539 121
rect 436 118 539 119
rect 614 121 677 122
rect 614 119 615 121
rect 617 119 674 121
rect 676 119 677 121
rect 614 118 677 119
rect 703 121 806 122
rect 703 119 704 121
rect 706 119 802 121
rect 804 119 806 121
rect 703 118 806 119
rect 881 121 944 122
rect 881 119 882 121
rect 884 119 941 121
rect 943 119 944 121
rect 881 118 944 119
rect 970 121 1073 122
rect 970 119 971 121
rect 973 119 1069 121
rect 1071 119 1073 121
rect 970 118 1073 119
rect 1148 121 1211 122
rect 1148 119 1149 121
rect 1151 119 1208 121
rect 1210 119 1211 121
rect 1148 118 1211 119
rect 1237 121 1340 122
rect 1237 119 1238 121
rect 1240 119 1336 121
rect 1338 119 1340 121
rect 1237 118 1340 119
rect 1415 121 1478 122
rect 1415 119 1416 121
rect 1418 119 1475 121
rect 1477 119 1478 121
rect 1415 118 1478 119
rect 1504 121 1607 122
rect 1504 119 1505 121
rect 1507 119 1603 121
rect 1605 119 1607 121
rect 1504 118 1607 119
rect 1682 121 1745 122
rect 1682 119 1683 121
rect 1685 119 1742 121
rect 1744 119 1745 121
rect 1682 118 1745 119
rect 1771 121 1874 122
rect 1771 119 1772 121
rect 1774 119 1870 121
rect 1872 119 1874 121
rect 1771 118 1874 119
rect 2057 121 2160 122
rect 2057 119 2058 121
rect 2060 119 2156 121
rect 2158 119 2160 121
rect 2057 118 2160 119
rect 299 117 307 118
rect 566 117 574 118
rect 833 117 841 118
rect 1100 117 1108 118
rect 1367 117 1375 118
rect 1634 117 1642 118
rect 1901 117 1909 118
rect 44 116 60 117
rect 44 114 45 116
rect 47 114 57 116
rect 59 114 60 116
rect 299 115 300 117
rect 302 115 304 117
rect 306 115 307 117
rect 299 114 307 115
rect 311 116 327 117
rect 311 114 312 116
rect 314 114 324 116
rect 326 114 327 116
rect 566 115 567 117
rect 569 115 571 117
rect 573 115 574 117
rect 566 114 574 115
rect 578 116 594 117
rect 578 114 579 116
rect 581 114 591 116
rect 593 114 594 116
rect 833 115 834 117
rect 836 115 838 117
rect 840 115 841 117
rect 833 114 841 115
rect 845 116 861 117
rect 845 114 846 116
rect 848 114 858 116
rect 860 114 861 116
rect 1100 115 1101 117
rect 1103 115 1105 117
rect 1107 115 1108 117
rect 1100 114 1108 115
rect 1112 116 1128 117
rect 1112 114 1113 116
rect 1115 114 1125 116
rect 1127 114 1128 116
rect 1367 115 1368 117
rect 1370 115 1372 117
rect 1374 115 1375 117
rect 1367 114 1375 115
rect 1379 116 1395 117
rect 1379 114 1380 116
rect 1382 114 1392 116
rect 1394 114 1395 116
rect 1634 115 1635 117
rect 1637 115 1639 117
rect 1641 115 1642 117
rect 1634 114 1642 115
rect 1646 116 1662 117
rect 1646 114 1647 116
rect 1649 114 1659 116
rect 1661 114 1662 116
rect 1901 115 1902 117
rect 1904 115 1906 117
rect 1908 115 1909 117
rect 1901 114 1909 115
rect 2187 117 2195 118
rect 2187 115 2188 117
rect 2190 115 2192 117
rect 2194 115 2195 117
rect 2187 114 2195 115
rect 44 113 60 114
rect 88 113 214 114
rect 311 113 327 114
rect 355 113 481 114
rect 578 113 594 114
rect 622 113 748 114
rect 845 113 861 114
rect 889 113 1015 114
rect 1112 113 1128 114
rect 1156 113 1282 114
rect 1379 113 1395 114
rect 1423 113 1549 114
rect 1646 113 1662 114
rect 1690 113 1816 114
rect 88 111 89 113
rect 91 111 211 113
rect 213 111 214 113
rect 88 110 214 111
rect 355 111 356 113
rect 358 111 478 113
rect 480 111 481 113
rect 355 110 481 111
rect 622 111 623 113
rect 625 111 745 113
rect 747 111 748 113
rect 622 110 748 111
rect 889 111 890 113
rect 892 111 1012 113
rect 1014 111 1015 113
rect 889 110 1015 111
rect 1156 111 1157 113
rect 1159 111 1279 113
rect 1281 111 1282 113
rect 1156 110 1282 111
rect 1423 111 1424 113
rect 1426 111 1546 113
rect 1548 111 1549 113
rect 1423 110 1549 111
rect 1690 111 1691 113
rect 1693 111 1813 113
rect 1815 111 1816 113
rect 1690 110 1816 111
rect 1860 113 1876 114
rect 1976 113 2102 114
rect 1860 111 1861 113
rect 1863 111 1873 113
rect 1875 111 1876 113
rect 1860 110 1876 111
rect 1924 112 1932 113
rect 1924 110 1925 112
rect 1927 110 1929 112
rect 1931 110 1932 112
rect 1976 111 1977 113
rect 1979 111 2099 113
rect 2101 111 2102 113
rect 2206 113 2210 114
rect 1976 110 2102 111
rect 2146 111 2150 112
rect 1924 109 1932 110
rect 2146 109 2147 111
rect 2149 110 2150 111
rect 2206 111 2207 113
rect 2209 111 2210 113
rect 2206 110 2210 111
rect 2149 109 2210 110
rect 2146 106 2210 109
rect 2275 113 2279 114
rect 2275 111 2276 113
rect 2278 111 2279 113
rect 260 104 339 105
rect 260 102 261 104
rect 263 102 336 104
rect 338 102 339 104
rect 260 101 339 102
rect 527 104 606 105
rect 527 102 528 104
rect 530 102 603 104
rect 605 102 606 104
rect 527 101 606 102
rect 794 104 873 105
rect 794 102 795 104
rect 797 102 870 104
rect 872 102 873 104
rect 794 101 873 102
rect 1061 104 1140 105
rect 1061 102 1062 104
rect 1064 102 1137 104
rect 1139 102 1140 104
rect 1061 101 1140 102
rect 1328 104 1407 105
rect 1328 102 1329 104
rect 1331 102 1404 104
rect 1406 102 1407 104
rect 1328 101 1407 102
rect 1595 104 1674 105
rect 1595 102 1596 104
rect 1598 102 1671 104
rect 1673 102 1674 104
rect 1595 101 1674 102
rect 2275 89 2279 111
rect 2275 87 2276 89
rect 2278 87 2279 89
rect 1862 79 1868 80
rect 1862 77 1865 79
rect 1867 77 1868 79
rect 260 74 355 75
rect 260 72 261 74
rect 263 72 352 74
rect 354 72 355 74
rect 260 71 355 72
rect 527 74 622 75
rect 527 72 528 74
rect 530 72 619 74
rect 621 72 622 74
rect 527 71 622 72
rect 794 74 889 75
rect 794 72 795 74
rect 797 72 886 74
rect 888 72 889 74
rect 794 71 889 72
rect 1061 74 1156 75
rect 1061 72 1062 74
rect 1064 72 1153 74
rect 1155 72 1156 74
rect 1061 71 1156 72
rect 1328 74 1423 75
rect 1328 72 1329 74
rect 1331 72 1420 74
rect 1422 72 1423 74
rect 1328 71 1423 72
rect 1595 74 1690 75
rect 1595 72 1596 74
rect 1598 72 1687 74
rect 1689 72 1690 74
rect 1595 71 1690 72
rect 1862 74 1868 77
rect 1862 72 1863 74
rect 1865 72 1868 74
rect 1862 71 1868 72
rect 2148 74 2213 75
rect 2148 72 2149 74
rect 2151 72 2213 74
rect 2148 71 2213 72
rect 1924 66 1932 67
rect 88 65 214 66
rect 88 63 89 65
rect 91 63 211 65
rect 213 63 214 65
rect 355 65 481 66
rect 88 62 214 63
rect 218 63 271 64
rect 2 61 20 62
rect 2 59 3 61
rect 5 59 17 61
rect 19 59 20 61
rect 2 58 20 59
rect 218 61 268 63
rect 270 61 271 63
rect 355 63 356 65
rect 358 63 478 65
rect 480 63 481 65
rect 622 65 748 66
rect 355 62 481 63
rect 485 63 538 64
rect 218 60 271 61
rect 485 61 535 63
rect 537 61 538 63
rect 622 63 623 65
rect 625 63 745 65
rect 747 63 748 65
rect 889 65 1015 66
rect 622 62 748 63
rect 752 63 805 64
rect 485 60 538 61
rect 752 61 802 63
rect 804 61 805 63
rect 889 63 890 65
rect 892 63 1012 65
rect 1014 63 1015 65
rect 1156 65 1282 66
rect 889 62 1015 63
rect 1019 63 1072 64
rect 752 60 805 61
rect 1019 61 1069 63
rect 1071 61 1072 63
rect 1156 63 1157 65
rect 1159 63 1279 65
rect 1281 63 1282 65
rect 1423 65 1549 66
rect 1156 62 1282 63
rect 1286 63 1339 64
rect 1019 60 1072 61
rect 1286 61 1336 63
rect 1338 61 1339 63
rect 1423 63 1424 65
rect 1426 63 1546 65
rect 1548 63 1549 65
rect 1690 65 1816 66
rect 1423 62 1549 63
rect 1553 63 1606 64
rect 1286 60 1339 61
rect 1553 61 1603 63
rect 1605 61 1606 63
rect 1690 63 1691 65
rect 1693 63 1813 65
rect 1815 63 1816 65
rect 1924 64 1925 66
rect 1927 64 1929 66
rect 1931 64 1932 66
rect 1690 62 1816 63
rect 1820 63 1873 64
rect 1924 63 1932 64
rect 1976 65 2102 66
rect 1976 63 1977 65
rect 1979 63 2099 65
rect 2101 63 2102 65
rect 2209 65 2213 71
rect 1553 60 1606 61
rect 1820 61 1870 63
rect 1872 61 1873 63
rect 1976 62 2102 63
rect 2106 63 2159 64
rect 1820 60 1873 61
rect 2106 61 2156 63
rect 2158 61 2159 63
rect 2209 63 2210 65
rect 2212 63 2213 65
rect 2209 62 2213 63
rect 2275 65 2279 87
rect 2310 85 2318 86
rect 2310 83 2311 85
rect 2313 83 2315 85
rect 2317 83 2318 85
rect 2310 82 2318 83
rect 2275 63 2276 65
rect 2278 63 2279 65
rect 2275 62 2279 63
rect 2106 60 2159 61
rect 218 58 222 60
rect 485 58 489 60
rect 752 58 756 60
rect 1019 58 1023 60
rect 1286 58 1290 60
rect 1553 58 1557 60
rect 1820 58 1824 60
rect 2106 58 2110 60
rect 80 57 142 58
rect 80 55 81 57
rect 83 55 139 57
rect 141 55 142 57
rect 80 54 142 55
rect 169 57 222 58
rect 169 55 170 57
rect 172 55 222 57
rect 169 54 222 55
rect 347 57 409 58
rect 347 55 348 57
rect 350 55 406 57
rect 408 55 409 57
rect 347 54 409 55
rect 436 57 489 58
rect 436 55 437 57
rect 439 55 489 57
rect 436 54 489 55
rect 614 57 676 58
rect 614 55 615 57
rect 617 55 673 57
rect 675 55 676 57
rect 614 54 676 55
rect 703 57 756 58
rect 703 55 704 57
rect 706 55 756 57
rect 703 54 756 55
rect 881 57 943 58
rect 881 55 882 57
rect 884 55 940 57
rect 942 55 943 57
rect 881 54 943 55
rect 970 57 1023 58
rect 970 55 971 57
rect 973 55 1023 57
rect 970 54 1023 55
rect 1148 57 1210 58
rect 1148 55 1149 57
rect 1151 55 1207 57
rect 1209 55 1210 57
rect 1148 54 1210 55
rect 1237 57 1290 58
rect 1237 55 1238 57
rect 1240 55 1290 57
rect 1237 54 1290 55
rect 1415 57 1477 58
rect 1415 55 1416 57
rect 1418 55 1474 57
rect 1476 55 1477 57
rect 1415 54 1477 55
rect 1504 57 1557 58
rect 1504 55 1505 57
rect 1507 55 1557 57
rect 1504 54 1557 55
rect 1682 57 1744 58
rect 1682 55 1683 57
rect 1685 55 1741 57
rect 1743 55 1744 57
rect 1682 54 1744 55
rect 1771 57 1824 58
rect 1771 55 1772 57
rect 1774 55 1824 57
rect 1771 54 1824 55
rect 2057 57 2110 58
rect 2057 55 2058 57
rect 2060 55 2110 57
rect 2057 54 2110 55
rect 227 52 307 53
rect 227 50 228 52
rect 230 50 304 52
rect 306 50 307 52
rect 494 52 574 53
rect 494 50 495 52
rect 497 50 571 52
rect 573 50 574 52
rect 761 52 841 53
rect 761 50 762 52
rect 764 50 838 52
rect 840 50 841 52
rect 1028 52 1108 53
rect 1028 50 1029 52
rect 1031 50 1105 52
rect 1107 50 1108 52
rect 1295 52 1375 53
rect 1295 50 1296 52
rect 1298 50 1372 52
rect 1374 50 1375 52
rect 1562 52 1642 53
rect 1562 50 1563 52
rect 1565 50 1639 52
rect 1641 50 1642 52
rect 1829 52 1909 53
rect 1829 50 1830 52
rect 1832 50 1906 52
rect 1908 50 1909 52
rect 2115 52 2195 53
rect 2115 50 2116 52
rect 2118 50 2192 52
rect 2194 50 2195 52
rect 40 49 136 50
rect 227 49 307 50
rect 335 49 403 50
rect 494 49 574 50
rect 602 49 670 50
rect 761 49 841 50
rect 869 49 937 50
rect 1028 49 1108 50
rect 1136 49 1204 50
rect 1295 49 1375 50
rect 1403 49 1471 50
rect 1562 49 1642 50
rect 1670 49 1738 50
rect 1829 49 1909 50
rect 1968 49 2021 50
rect 2115 49 2195 50
rect 2219 50 2239 51
rect 40 47 41 49
rect 43 47 133 49
rect 135 47 136 49
rect 40 46 136 47
rect 335 47 336 49
rect 338 47 400 49
rect 402 47 403 49
rect 335 46 403 47
rect 602 47 603 49
rect 605 47 667 49
rect 669 47 670 49
rect 602 46 670 47
rect 869 47 870 49
rect 872 47 934 49
rect 936 47 937 49
rect 869 46 937 47
rect 1136 47 1137 49
rect 1139 47 1201 49
rect 1203 47 1204 49
rect 1136 46 1204 47
rect 1403 47 1404 49
rect 1406 47 1468 49
rect 1470 47 1471 49
rect 1403 46 1471 47
rect 1670 47 1671 49
rect 1673 47 1735 49
rect 1737 47 1738 49
rect 1670 46 1738 47
rect 1968 47 1969 49
rect 1971 47 2018 49
rect 2020 47 2021 49
rect 2219 48 2220 50
rect 2222 48 2236 50
rect 2238 48 2239 50
rect 2219 47 2239 48
rect 2299 50 2307 51
rect 2299 48 2300 50
rect 2302 48 2304 50
rect 2306 48 2307 50
rect 2299 47 2307 48
rect 1968 46 2021 47
rect 179 44 271 45
rect 179 42 180 44
rect 182 42 268 44
rect 270 42 271 44
rect 446 44 538 45
rect 446 42 447 44
rect 449 42 535 44
rect 537 42 538 44
rect 713 44 805 45
rect 713 42 714 44
rect 716 42 802 44
rect 804 42 805 44
rect 980 44 1072 45
rect 980 42 981 44
rect 983 42 1069 44
rect 1071 42 1072 44
rect 1247 44 1339 45
rect 1247 42 1248 44
rect 1250 42 1336 44
rect 1338 42 1339 44
rect 1514 44 1606 45
rect 1514 42 1515 44
rect 1517 42 1603 44
rect 1605 42 1606 44
rect 1781 44 1873 45
rect 1781 42 1782 44
rect 1784 42 1870 44
rect 1872 42 1873 44
rect 44 41 52 42
rect 179 41 271 42
rect 311 41 319 42
rect 446 41 538 42
rect 578 41 586 42
rect 713 41 805 42
rect 845 41 853 42
rect 980 41 1072 42
rect 1112 41 1120 42
rect 1247 41 1339 42
rect 1379 41 1387 42
rect 1514 41 1606 42
rect 1646 41 1654 42
rect 1781 41 1873 42
rect 2067 44 2159 45
rect 2067 42 2068 44
rect 2070 42 2156 44
rect 2158 42 2159 44
rect 2067 41 2159 42
rect 44 39 45 41
rect 47 39 49 41
rect 51 39 52 41
rect 44 38 52 39
rect 311 39 312 41
rect 314 39 316 41
rect 318 39 319 41
rect 311 38 319 39
rect 578 39 579 41
rect 581 39 583 41
rect 585 39 586 41
rect 578 38 586 39
rect 845 39 846 41
rect 848 39 850 41
rect 852 39 853 41
rect 845 38 853 39
rect 1112 39 1113 41
rect 1115 39 1117 41
rect 1119 39 1120 41
rect 1112 38 1120 39
rect 1379 39 1380 41
rect 1382 39 1384 41
rect 1386 39 1387 41
rect 1379 38 1387 39
rect 1646 39 1647 41
rect 1649 39 1651 41
rect 1653 39 1654 41
rect 1646 38 1654 39
rect 290 33 294 34
rect 290 31 291 33
rect 293 31 294 33
rect 183 -6 271 -5
rect 183 -8 268 -6
rect 270 -8 271 -6
rect 183 -9 271 -8
rect 179 -10 187 -9
rect 2 -12 12 -11
rect 2 -14 3 -12
rect 5 -14 9 -12
rect 11 -14 12 -12
rect 179 -12 180 -10
rect 182 -12 187 -10
rect 179 -13 187 -12
rect 290 -14 294 31
rect 557 33 561 34
rect 557 31 558 33
rect 560 31 561 33
rect 450 -6 538 -5
rect 450 -8 535 -6
rect 537 -8 538 -6
rect 450 -9 538 -8
rect 446 -10 454 -9
rect 446 -12 447 -10
rect 449 -12 454 -10
rect 446 -13 454 -12
rect 557 -14 561 31
rect 824 33 828 34
rect 824 31 825 33
rect 827 31 828 33
rect 717 -6 805 -5
rect 717 -8 802 -6
rect 804 -8 805 -6
rect 717 -9 805 -8
rect 713 -10 721 -9
rect 713 -12 714 -10
rect 716 -12 721 -10
rect 713 -13 721 -12
rect 824 -14 828 31
rect 1091 33 1095 34
rect 1091 31 1092 33
rect 1094 31 1095 33
rect 984 -6 1072 -5
rect 984 -8 1069 -6
rect 1071 -8 1072 -6
rect 984 -9 1072 -8
rect 980 -10 988 -9
rect 980 -12 981 -10
rect 983 -12 988 -10
rect 980 -13 988 -12
rect 1091 -14 1095 31
rect 1358 33 1362 34
rect 1358 31 1359 33
rect 1361 31 1362 33
rect 1251 -6 1339 -5
rect 1251 -8 1336 -6
rect 1338 -8 1339 -6
rect 1251 -9 1339 -8
rect 1247 -10 1255 -9
rect 1247 -12 1248 -10
rect 1250 -12 1255 -10
rect 1247 -13 1255 -12
rect 1358 -14 1362 31
rect 1625 33 1629 34
rect 1625 31 1626 33
rect 1628 31 1629 33
rect 1518 -6 1606 -5
rect 1518 -8 1603 -6
rect 1605 -8 1606 -6
rect 1518 -9 1606 -8
rect 1514 -10 1522 -9
rect 1514 -12 1515 -10
rect 1517 -12 1522 -10
rect 1514 -13 1522 -12
rect 1625 -14 1629 31
rect 1892 33 1896 34
rect 1892 31 1893 33
rect 1895 31 1896 33
rect 1785 -6 1873 -5
rect 1785 -8 1870 -6
rect 1872 -8 1873 -6
rect 1785 -9 1873 -8
rect 1781 -10 1789 -9
rect 1781 -12 1782 -10
rect 1784 -12 1789 -10
rect 1781 -13 1789 -12
rect 1892 -14 1896 31
rect 2179 33 2183 34
rect 2179 31 2180 33
rect 2182 31 2183 33
rect 2105 -6 2159 -5
rect 2105 -8 2156 -6
rect 2158 -8 2159 -6
rect 2105 -9 2159 -8
rect 2067 -10 2111 -9
rect 2067 -12 2068 -10
rect 2070 -12 2111 -10
rect 2067 -13 2111 -12
rect 2179 -14 2183 31
rect 2319 23 2327 24
rect 2319 21 2320 23
rect 2322 21 2324 23
rect 2326 21 2327 23
rect 2319 20 2327 21
rect 2 -15 12 -14
rect 45 -15 124 -14
rect 45 -17 121 -15
rect 123 -17 124 -15
rect 40 -18 124 -17
rect 226 -15 295 -14
rect 226 -17 227 -15
rect 229 -17 295 -15
rect 226 -18 295 -17
rect 351 -15 391 -14
rect 351 -17 352 -15
rect 354 -17 388 -15
rect 390 -17 391 -15
rect 351 -18 391 -17
rect 493 -15 562 -14
rect 493 -17 494 -15
rect 496 -17 562 -15
rect 493 -18 562 -17
rect 618 -15 658 -14
rect 618 -17 619 -15
rect 621 -17 655 -15
rect 657 -17 658 -15
rect 618 -18 658 -17
rect 760 -15 829 -14
rect 760 -17 761 -15
rect 763 -17 829 -15
rect 760 -18 829 -17
rect 885 -15 925 -14
rect 885 -17 886 -15
rect 888 -17 922 -15
rect 924 -17 925 -15
rect 885 -18 925 -17
rect 1027 -15 1096 -14
rect 1027 -17 1028 -15
rect 1030 -17 1096 -15
rect 1027 -18 1096 -17
rect 1152 -15 1192 -14
rect 1152 -17 1153 -15
rect 1155 -17 1189 -15
rect 1191 -17 1192 -15
rect 1152 -18 1192 -17
rect 1294 -15 1363 -14
rect 1294 -17 1295 -15
rect 1297 -17 1363 -15
rect 1294 -18 1363 -17
rect 1419 -15 1459 -14
rect 1419 -17 1420 -15
rect 1422 -17 1456 -15
rect 1458 -17 1459 -15
rect 1419 -18 1459 -17
rect 1561 -15 1630 -14
rect 1561 -17 1562 -15
rect 1564 -17 1630 -15
rect 1561 -18 1630 -17
rect 1686 -15 1726 -14
rect 1686 -17 1687 -15
rect 1689 -17 1723 -15
rect 1725 -17 1726 -15
rect 1686 -18 1726 -17
rect 1828 -15 1897 -14
rect 1828 -17 1829 -15
rect 1831 -17 1897 -15
rect 1828 -18 1897 -17
rect 1968 -15 2021 -14
rect 1968 -17 1969 -15
rect 1971 -17 2018 -15
rect 2020 -17 2021 -15
rect 1968 -18 2021 -17
rect 2115 -15 2183 -14
rect 2115 -17 2116 -15
rect 2118 -17 2183 -15
rect 2235 -14 2239 -13
rect 2235 -16 2236 -14
rect 2238 -16 2239 -14
rect 2115 -18 2183 -17
rect 2227 -17 2239 -16
rect 2299 -14 2307 -13
rect 2299 -16 2300 -14
rect 2302 -16 2304 -14
rect 2306 -16 2307 -14
rect 2299 -17 2307 -16
rect 40 -20 41 -18
rect 43 -20 49 -18
rect 2227 -19 2228 -17
rect 2230 -19 2239 -17
rect 2227 -20 2239 -19
rect 40 -21 49 -20
rect 80 -23 142 -22
rect 80 -25 81 -23
rect 83 -25 139 -23
rect 141 -25 142 -23
rect 80 -26 142 -25
rect 169 -23 272 -22
rect 169 -25 170 -23
rect 172 -25 268 -23
rect 270 -25 272 -23
rect 169 -26 272 -25
rect 347 -23 409 -22
rect 347 -25 348 -23
rect 350 -25 406 -23
rect 408 -25 409 -23
rect 347 -26 409 -25
rect 436 -23 539 -22
rect 436 -25 437 -23
rect 439 -25 535 -23
rect 537 -25 539 -23
rect 436 -26 539 -25
rect 614 -23 676 -22
rect 614 -25 615 -23
rect 617 -25 673 -23
rect 675 -25 676 -23
rect 614 -26 676 -25
rect 703 -23 806 -22
rect 703 -25 704 -23
rect 706 -25 802 -23
rect 804 -25 806 -23
rect 703 -26 806 -25
rect 881 -23 943 -22
rect 881 -25 882 -23
rect 884 -25 940 -23
rect 942 -25 943 -23
rect 881 -26 943 -25
rect 970 -23 1073 -22
rect 970 -25 971 -23
rect 973 -25 1069 -23
rect 1071 -25 1073 -23
rect 970 -26 1073 -25
rect 1148 -23 1210 -22
rect 1148 -25 1149 -23
rect 1151 -25 1207 -23
rect 1209 -25 1210 -23
rect 1148 -26 1210 -25
rect 1237 -23 1340 -22
rect 1237 -25 1238 -23
rect 1240 -25 1336 -23
rect 1338 -25 1340 -23
rect 1237 -26 1340 -25
rect 1415 -23 1477 -22
rect 1415 -25 1416 -23
rect 1418 -25 1474 -23
rect 1476 -25 1477 -23
rect 1415 -26 1477 -25
rect 1504 -23 1607 -22
rect 1504 -25 1505 -23
rect 1507 -25 1603 -23
rect 1605 -25 1607 -23
rect 1504 -26 1607 -25
rect 1682 -23 1744 -22
rect 1682 -25 1683 -23
rect 1685 -25 1741 -23
rect 1743 -25 1744 -23
rect 1682 -26 1744 -25
rect 1771 -23 1874 -22
rect 1771 -25 1772 -23
rect 1774 -25 1870 -23
rect 1872 -25 1874 -23
rect 1771 -26 1874 -25
rect 2057 -23 2160 -22
rect 2057 -25 2058 -23
rect 2060 -25 2156 -23
rect 2158 -25 2160 -23
rect 2057 -26 2160 -25
rect 299 -27 307 -26
rect 44 -29 60 -28
rect 44 -31 45 -29
rect 47 -31 57 -29
rect 59 -31 60 -29
rect 299 -29 300 -27
rect 302 -29 304 -27
rect 306 -29 307 -27
rect 566 -27 574 -26
rect 299 -30 307 -29
rect 311 -29 327 -28
rect 44 -33 60 -31
rect 88 -31 214 -30
rect 88 -33 89 -31
rect 91 -33 211 -31
rect 213 -33 214 -31
rect 88 -34 214 -33
rect 258 -31 262 -30
rect 258 -33 259 -31
rect 261 -33 262 -31
rect 311 -31 312 -29
rect 314 -31 324 -29
rect 326 -31 327 -29
rect 566 -29 567 -27
rect 569 -29 571 -27
rect 573 -29 574 -27
rect 833 -27 841 -26
rect 566 -30 574 -29
rect 578 -29 594 -28
rect 311 -33 327 -31
rect 355 -31 481 -30
rect 355 -33 356 -31
rect 358 -33 478 -31
rect 480 -33 481 -31
rect 258 -39 262 -33
rect 355 -34 481 -33
rect 525 -31 529 -30
rect 525 -33 526 -31
rect 528 -33 529 -31
rect 578 -31 579 -29
rect 581 -31 591 -29
rect 593 -31 594 -29
rect 833 -29 834 -27
rect 836 -29 838 -27
rect 840 -29 841 -27
rect 1100 -27 1108 -26
rect 833 -30 841 -29
rect 845 -29 861 -28
rect 578 -33 594 -31
rect 622 -31 748 -30
rect 622 -33 623 -31
rect 625 -33 745 -31
rect 747 -33 748 -31
rect 525 -39 529 -33
rect 622 -34 748 -33
rect 792 -31 796 -30
rect 792 -33 793 -31
rect 795 -33 796 -31
rect 845 -31 846 -29
rect 848 -31 858 -29
rect 860 -31 861 -29
rect 1100 -29 1101 -27
rect 1103 -29 1105 -27
rect 1107 -29 1108 -27
rect 1367 -27 1375 -26
rect 1100 -30 1108 -29
rect 1112 -29 1128 -28
rect 845 -33 861 -31
rect 889 -31 1015 -30
rect 889 -33 890 -31
rect 892 -33 1012 -31
rect 1014 -33 1015 -31
rect 792 -39 796 -33
rect 889 -34 1015 -33
rect 1059 -31 1063 -30
rect 1059 -33 1060 -31
rect 1062 -33 1063 -31
rect 1112 -31 1113 -29
rect 1115 -31 1125 -29
rect 1127 -31 1128 -29
rect 1367 -29 1368 -27
rect 1370 -29 1372 -27
rect 1374 -29 1375 -27
rect 1634 -27 1642 -26
rect 1367 -30 1375 -29
rect 1379 -29 1395 -28
rect 1112 -33 1128 -31
rect 1156 -31 1282 -30
rect 1156 -33 1157 -31
rect 1159 -33 1279 -31
rect 1281 -33 1282 -31
rect 1059 -39 1063 -33
rect 1156 -34 1282 -33
rect 1326 -31 1330 -30
rect 1326 -33 1327 -31
rect 1329 -33 1330 -31
rect 1379 -31 1380 -29
rect 1382 -31 1392 -29
rect 1394 -31 1395 -29
rect 1634 -29 1635 -27
rect 1637 -29 1639 -27
rect 1641 -29 1642 -27
rect 1901 -27 1909 -26
rect 1634 -30 1642 -29
rect 1646 -29 1662 -28
rect 1379 -33 1395 -31
rect 1423 -31 1549 -30
rect 1423 -33 1424 -31
rect 1426 -33 1546 -31
rect 1548 -33 1549 -31
rect 1326 -39 1330 -33
rect 1423 -34 1549 -33
rect 1593 -31 1597 -30
rect 1593 -33 1594 -31
rect 1596 -33 1597 -31
rect 1646 -31 1647 -29
rect 1649 -31 1659 -29
rect 1661 -31 1662 -29
rect 1901 -29 1902 -27
rect 1904 -29 1906 -27
rect 1908 -29 1909 -27
rect 1901 -30 1909 -29
rect 2187 -27 2195 -26
rect 2187 -29 2188 -27
rect 2190 -29 2192 -27
rect 2194 -29 2195 -27
rect 2187 -30 2195 -29
rect 1646 -33 1662 -31
rect 1690 -31 1816 -30
rect 1976 -31 2102 -30
rect 1690 -33 1691 -31
rect 1693 -33 1813 -31
rect 1815 -33 1816 -31
rect 1593 -39 1597 -33
rect 1690 -34 1816 -33
rect 1856 -32 1864 -31
rect 1856 -34 1857 -32
rect 1859 -34 1861 -32
rect 1863 -34 1864 -32
rect 1856 -35 1864 -34
rect 1924 -32 1932 -31
rect 1924 -34 1925 -32
rect 1927 -34 1929 -32
rect 1931 -34 1932 -32
rect 1976 -33 1977 -31
rect 1979 -33 2099 -31
rect 2101 -33 2102 -31
rect 1976 -34 2102 -33
rect 2146 -31 2150 -30
rect 2146 -33 2147 -31
rect 2149 -33 2150 -31
rect 2146 -34 2150 -33
rect 2209 -31 2213 -30
rect 2209 -33 2210 -31
rect 2212 -33 2213 -31
rect 2209 -34 2213 -33
rect 1924 -35 1932 -34
rect 2146 -38 2213 -34
rect 2275 -31 2279 -30
rect 2275 -33 2276 -31
rect 2278 -33 2279 -31
rect 258 -40 339 -39
rect 258 -42 336 -40
rect 338 -42 339 -40
rect 258 -43 339 -42
rect 525 -40 606 -39
rect 525 -42 603 -40
rect 605 -42 606 -40
rect 525 -43 606 -42
rect 792 -40 873 -39
rect 792 -42 870 -40
rect 872 -42 873 -40
rect 792 -43 873 -42
rect 1059 -40 1140 -39
rect 1059 -42 1137 -40
rect 1139 -42 1140 -40
rect 1059 -43 1140 -42
rect 1326 -40 1407 -39
rect 1326 -42 1404 -40
rect 1406 -42 1407 -40
rect 1326 -43 1407 -42
rect 1593 -40 1674 -39
rect 1593 -42 1671 -40
rect 1673 -42 1674 -40
rect 1593 -43 1674 -42
rect 2275 -55 2279 -33
rect 2275 -57 2276 -55
rect 2278 -57 2279 -55
rect 260 -70 355 -69
rect 260 -72 261 -70
rect 263 -72 352 -70
rect 354 -72 355 -70
rect 260 -73 355 -72
rect 527 -70 622 -69
rect 527 -72 528 -70
rect 530 -72 619 -70
rect 621 -72 622 -70
rect 527 -73 622 -72
rect 794 -70 889 -69
rect 794 -72 795 -70
rect 797 -72 886 -70
rect 888 -72 889 -70
rect 794 -73 889 -72
rect 1061 -70 1156 -69
rect 1061 -72 1062 -70
rect 1064 -72 1153 -70
rect 1155 -72 1156 -70
rect 1061 -73 1156 -72
rect 1328 -70 1423 -69
rect 1328 -72 1329 -70
rect 1331 -72 1420 -70
rect 1422 -72 1423 -70
rect 1328 -73 1423 -72
rect 1595 -70 1690 -69
rect 1595 -72 1596 -70
rect 1598 -72 1687 -70
rect 1689 -72 1690 -70
rect 1595 -73 1690 -72
rect 1848 -70 1866 -69
rect 1848 -72 1849 -70
rect 1851 -72 1863 -70
rect 1865 -72 1866 -70
rect 1848 -73 1866 -72
rect 2148 -70 2213 -69
rect 2148 -72 2149 -70
rect 2151 -72 2213 -70
rect 2148 -73 2213 -72
rect 1924 -78 1932 -77
rect 88 -79 214 -78
rect 88 -81 89 -79
rect 91 -81 211 -79
rect 213 -81 214 -79
rect 355 -79 481 -78
rect 88 -82 214 -81
rect 218 -81 271 -80
rect 2 -83 20 -82
rect 2 -85 3 -83
rect 5 -85 17 -83
rect 19 -85 20 -83
rect 2 -86 20 -85
rect 218 -83 268 -81
rect 270 -83 271 -81
rect 355 -81 356 -79
rect 358 -81 478 -79
rect 480 -81 481 -79
rect 622 -79 748 -78
rect 355 -82 481 -81
rect 485 -81 538 -80
rect 218 -84 271 -83
rect 485 -83 535 -81
rect 537 -83 538 -81
rect 622 -81 623 -79
rect 625 -81 745 -79
rect 747 -81 748 -79
rect 889 -79 1015 -78
rect 622 -82 748 -81
rect 752 -81 805 -80
rect 485 -84 538 -83
rect 752 -83 802 -81
rect 804 -83 805 -81
rect 889 -81 890 -79
rect 892 -81 1012 -79
rect 1014 -81 1015 -79
rect 1156 -79 1282 -78
rect 889 -82 1015 -81
rect 1019 -81 1072 -80
rect 752 -84 805 -83
rect 1019 -83 1069 -81
rect 1071 -83 1072 -81
rect 1156 -81 1157 -79
rect 1159 -81 1279 -79
rect 1281 -81 1282 -79
rect 1423 -79 1549 -78
rect 1156 -82 1282 -81
rect 1286 -81 1339 -80
rect 1019 -84 1072 -83
rect 1286 -83 1336 -81
rect 1338 -83 1339 -81
rect 1423 -81 1424 -79
rect 1426 -81 1546 -79
rect 1548 -81 1549 -79
rect 1690 -79 1816 -78
rect 1423 -82 1549 -81
rect 1553 -81 1606 -80
rect 1286 -84 1339 -83
rect 1553 -83 1603 -81
rect 1605 -83 1606 -81
rect 1690 -81 1691 -79
rect 1693 -81 1813 -79
rect 1815 -81 1816 -79
rect 1924 -80 1925 -78
rect 1927 -80 1929 -78
rect 1931 -80 1932 -78
rect 1690 -82 1816 -81
rect 1820 -81 1873 -80
rect 1924 -81 1932 -80
rect 1976 -79 2102 -78
rect 1976 -81 1977 -79
rect 1979 -81 2099 -79
rect 2101 -81 2102 -79
rect 2209 -79 2213 -73
rect 1553 -84 1606 -83
rect 1820 -83 1870 -81
rect 1872 -83 1873 -81
rect 1976 -82 2102 -81
rect 2106 -81 2159 -80
rect 1820 -84 1873 -83
rect 2106 -83 2156 -81
rect 2158 -83 2159 -81
rect 2209 -81 2210 -79
rect 2212 -81 2213 -79
rect 2209 -82 2213 -81
rect 2275 -79 2279 -57
rect 2310 -59 2318 -58
rect 2310 -61 2311 -59
rect 2313 -61 2315 -59
rect 2317 -61 2318 -59
rect 2310 -62 2318 -61
rect 2275 -81 2276 -79
rect 2278 -81 2279 -79
rect 2275 -82 2279 -81
rect 2106 -84 2159 -83
rect 218 -86 222 -84
rect 485 -86 489 -84
rect 752 -86 756 -84
rect 1019 -86 1023 -84
rect 1286 -86 1290 -84
rect 1553 -86 1557 -84
rect 1820 -86 1824 -84
rect 2106 -86 2110 -84
rect 80 -87 142 -86
rect 80 -89 81 -87
rect 83 -89 139 -87
rect 141 -89 142 -87
rect 80 -90 142 -89
rect 169 -87 222 -86
rect 169 -89 170 -87
rect 172 -89 222 -87
rect 169 -90 222 -89
rect 347 -87 409 -86
rect 347 -89 348 -87
rect 350 -89 406 -87
rect 408 -89 409 -87
rect 347 -90 409 -89
rect 436 -87 489 -86
rect 436 -89 437 -87
rect 439 -89 489 -87
rect 436 -90 489 -89
rect 614 -87 676 -86
rect 614 -89 615 -87
rect 617 -89 673 -87
rect 675 -89 676 -87
rect 614 -90 676 -89
rect 703 -87 756 -86
rect 703 -89 704 -87
rect 706 -89 756 -87
rect 703 -90 756 -89
rect 881 -87 943 -86
rect 881 -89 882 -87
rect 884 -89 940 -87
rect 942 -89 943 -87
rect 881 -90 943 -89
rect 970 -87 1023 -86
rect 970 -89 971 -87
rect 973 -89 1023 -87
rect 970 -90 1023 -89
rect 1148 -87 1210 -86
rect 1148 -89 1149 -87
rect 1151 -89 1207 -87
rect 1209 -89 1210 -87
rect 1148 -90 1210 -89
rect 1237 -87 1290 -86
rect 1237 -89 1238 -87
rect 1240 -89 1290 -87
rect 1237 -90 1290 -89
rect 1415 -87 1477 -86
rect 1415 -89 1416 -87
rect 1418 -89 1474 -87
rect 1476 -89 1477 -87
rect 1415 -90 1477 -89
rect 1504 -87 1557 -86
rect 1504 -89 1505 -87
rect 1507 -89 1557 -87
rect 1504 -90 1557 -89
rect 1682 -87 1744 -86
rect 1682 -89 1683 -87
rect 1685 -89 1741 -87
rect 1743 -89 1744 -87
rect 1682 -90 1744 -89
rect 1771 -87 1824 -86
rect 1771 -89 1772 -87
rect 1774 -89 1824 -87
rect 1771 -90 1824 -89
rect 2057 -87 2110 -86
rect 2057 -89 2058 -87
rect 2060 -89 2110 -87
rect 2057 -90 2110 -89
rect 227 -92 307 -91
rect 227 -94 228 -92
rect 230 -94 304 -92
rect 306 -94 307 -92
rect 494 -92 574 -91
rect 494 -94 495 -92
rect 497 -94 571 -92
rect 573 -94 574 -92
rect 761 -92 841 -91
rect 761 -94 762 -92
rect 764 -94 838 -92
rect 840 -94 841 -92
rect 1028 -92 1108 -91
rect 1028 -94 1029 -92
rect 1031 -94 1105 -92
rect 1107 -94 1108 -92
rect 1295 -92 1375 -91
rect 1295 -94 1296 -92
rect 1298 -94 1372 -92
rect 1374 -94 1375 -92
rect 1562 -92 1642 -91
rect 1562 -94 1563 -92
rect 1565 -94 1639 -92
rect 1641 -94 1642 -92
rect 1829 -92 1909 -91
rect 1829 -94 1830 -92
rect 1832 -94 1906 -92
rect 1908 -94 1909 -92
rect 2115 -92 2195 -91
rect 2115 -94 2116 -92
rect 2118 -94 2192 -92
rect 2194 -94 2195 -92
rect 40 -95 137 -94
rect 227 -95 307 -94
rect 311 -95 404 -94
rect 494 -95 574 -94
rect 578 -95 671 -94
rect 761 -95 841 -94
rect 845 -95 938 -94
rect 1028 -95 1108 -94
rect 1112 -95 1205 -94
rect 1295 -95 1375 -94
rect 1379 -95 1472 -94
rect 1562 -95 1642 -94
rect 1646 -95 1739 -94
rect 1829 -95 1909 -94
rect 1968 -95 2021 -94
rect 2115 -95 2195 -94
rect 2235 -94 2239 -93
rect 40 -97 41 -95
rect 43 -97 134 -95
rect 136 -97 137 -95
rect 40 -98 137 -97
rect 311 -97 336 -95
rect 338 -97 401 -95
rect 403 -97 404 -95
rect 311 -98 404 -97
rect 578 -97 603 -95
rect 605 -97 668 -95
rect 670 -97 671 -95
rect 578 -98 671 -97
rect 845 -97 870 -95
rect 872 -97 935 -95
rect 937 -97 938 -95
rect 845 -98 938 -97
rect 1112 -97 1137 -95
rect 1139 -97 1202 -95
rect 1204 -97 1205 -95
rect 1112 -98 1205 -97
rect 1379 -97 1404 -95
rect 1406 -97 1469 -95
rect 1471 -97 1472 -95
rect 1379 -98 1472 -97
rect 1646 -97 1671 -95
rect 1673 -97 1736 -95
rect 1738 -97 1739 -95
rect 1646 -98 1739 -97
rect 1968 -97 1969 -95
rect 1971 -97 2018 -95
rect 2020 -97 2021 -95
rect 1968 -98 2021 -97
rect 2235 -96 2236 -94
rect 2238 -96 2239 -94
rect 2235 -99 2239 -96
rect 2299 -94 2307 -93
rect 2299 -96 2300 -94
rect 2302 -96 2304 -94
rect 2306 -96 2307 -94
rect 2299 -97 2307 -96
rect 179 -100 271 -99
rect 179 -102 180 -100
rect 182 -102 268 -100
rect 270 -102 271 -100
rect 446 -100 538 -99
rect 446 -102 447 -100
rect 449 -102 535 -100
rect 537 -102 538 -100
rect 713 -100 805 -99
rect 713 -102 714 -100
rect 716 -102 802 -100
rect 804 -102 805 -100
rect 980 -100 1072 -99
rect 980 -102 981 -100
rect 983 -102 1069 -100
rect 1071 -102 1072 -100
rect 1247 -100 1339 -99
rect 1247 -102 1248 -100
rect 1250 -102 1336 -100
rect 1338 -102 1339 -100
rect 1514 -100 1606 -99
rect 1514 -102 1515 -100
rect 1517 -102 1603 -100
rect 1605 -102 1606 -100
rect 1781 -100 1873 -99
rect 1781 -102 1782 -100
rect 1784 -102 1870 -100
rect 1872 -102 1873 -100
rect 44 -103 52 -102
rect 179 -103 271 -102
rect 311 -103 319 -102
rect 446 -103 538 -102
rect 578 -103 586 -102
rect 713 -103 805 -102
rect 845 -103 853 -102
rect 980 -103 1072 -102
rect 1112 -103 1120 -102
rect 1247 -103 1339 -102
rect 1379 -103 1387 -102
rect 1514 -103 1606 -102
rect 1646 -103 1654 -102
rect 1781 -103 1873 -102
rect 2067 -100 2159 -99
rect 2067 -102 2068 -100
rect 2070 -102 2156 -100
rect 2158 -102 2159 -100
rect 2235 -101 2236 -99
rect 2238 -101 2239 -99
rect 2235 -102 2239 -101
rect 2067 -103 2159 -102
rect 44 -105 45 -103
rect 47 -105 49 -103
rect 51 -105 52 -103
rect 44 -106 52 -105
rect 311 -105 312 -103
rect 314 -105 316 -103
rect 318 -105 319 -103
rect 311 -106 319 -105
rect 578 -105 579 -103
rect 581 -105 583 -103
rect 585 -105 586 -103
rect 578 -106 586 -105
rect 845 -105 846 -103
rect 848 -105 850 -103
rect 852 -105 853 -103
rect 845 -106 853 -105
rect 1112 -105 1113 -103
rect 1115 -105 1117 -103
rect 1119 -105 1120 -103
rect 1112 -106 1120 -105
rect 1379 -105 1380 -103
rect 1382 -105 1384 -103
rect 1386 -105 1387 -103
rect 1379 -106 1387 -105
rect 1646 -105 1647 -103
rect 1649 -105 1651 -103
rect 1653 -105 1654 -103
rect 1646 -106 1654 -105
rect 291 -111 295 -110
rect 291 -113 292 -111
rect 294 -113 295 -111
rect 219 -150 271 -149
rect 219 -152 268 -150
rect 270 -152 271 -150
rect 219 -153 271 -152
rect 179 -154 223 -153
rect 2 -156 12 -155
rect 2 -158 3 -156
rect 5 -158 9 -156
rect 11 -158 12 -156
rect 179 -156 180 -154
rect 182 -156 223 -154
rect 179 -157 223 -156
rect 291 -158 295 -113
rect 558 -111 562 -110
rect 558 -113 559 -111
rect 561 -113 562 -111
rect 486 -150 538 -149
rect 486 -152 535 -150
rect 537 -152 538 -150
rect 486 -153 538 -152
rect 446 -154 490 -153
rect 446 -156 447 -154
rect 449 -156 490 -154
rect 446 -157 490 -156
rect 558 -158 562 -113
rect 825 -111 829 -110
rect 825 -113 826 -111
rect 828 -113 829 -111
rect 753 -150 805 -149
rect 753 -152 802 -150
rect 804 -152 805 -150
rect 753 -153 805 -152
rect 713 -154 757 -153
rect 713 -156 714 -154
rect 716 -156 757 -154
rect 713 -157 757 -156
rect 825 -158 829 -113
rect 1092 -111 1096 -110
rect 1092 -113 1093 -111
rect 1095 -113 1096 -111
rect 1020 -150 1072 -149
rect 1020 -152 1069 -150
rect 1071 -152 1072 -150
rect 1020 -153 1072 -152
rect 980 -154 1024 -153
rect 980 -156 981 -154
rect 983 -156 1024 -154
rect 980 -157 1024 -156
rect 1092 -158 1096 -113
rect 1359 -111 1363 -110
rect 1359 -113 1360 -111
rect 1362 -113 1363 -111
rect 1287 -150 1339 -149
rect 1287 -152 1336 -150
rect 1338 -152 1339 -150
rect 1287 -153 1339 -152
rect 1247 -154 1291 -153
rect 1247 -156 1248 -154
rect 1250 -156 1291 -154
rect 1247 -157 1291 -156
rect 1359 -158 1363 -113
rect 1626 -111 1630 -110
rect 1626 -113 1627 -111
rect 1629 -113 1630 -111
rect 1554 -150 1606 -149
rect 1554 -152 1603 -150
rect 1605 -152 1606 -150
rect 1554 -153 1606 -152
rect 1514 -154 1558 -153
rect 1514 -156 1515 -154
rect 1517 -156 1558 -154
rect 1514 -157 1558 -156
rect 1626 -158 1630 -113
rect 1893 -111 1897 -110
rect 1893 -113 1894 -111
rect 1896 -113 1897 -111
rect 1821 -150 1873 -149
rect 1821 -152 1870 -150
rect 1872 -152 1873 -150
rect 1821 -153 1873 -152
rect 1781 -154 1825 -153
rect 1781 -156 1782 -154
rect 1784 -156 1825 -154
rect 1781 -157 1825 -156
rect 1893 -158 1897 -113
rect 2179 -111 2183 -110
rect 2179 -113 2180 -111
rect 2182 -113 2183 -111
rect 2107 -150 2159 -149
rect 2107 -152 2156 -150
rect 2158 -152 2159 -150
rect 2107 -153 2159 -152
rect 2067 -154 2111 -153
rect 2067 -156 2068 -154
rect 2070 -156 2111 -154
rect 2067 -157 2111 -156
rect 2179 -158 2183 -113
rect 2319 -121 2327 -120
rect 2319 -123 2320 -121
rect 2322 -123 2324 -121
rect 2326 -123 2327 -121
rect 2319 -124 2327 -123
rect 2 -159 12 -158
rect 39 -159 141 -158
rect 39 -161 41 -159
rect 43 -161 138 -159
rect 140 -161 141 -159
rect 39 -162 141 -161
rect 227 -159 295 -158
rect 227 -161 228 -159
rect 230 -161 295 -159
rect 227 -162 295 -161
rect 351 -159 408 -158
rect 351 -161 352 -159
rect 354 -161 405 -159
rect 407 -161 408 -159
rect 351 -162 408 -161
rect 494 -159 562 -158
rect 494 -161 495 -159
rect 497 -161 562 -159
rect 494 -162 562 -161
rect 618 -159 675 -158
rect 618 -161 619 -159
rect 621 -161 672 -159
rect 674 -161 675 -159
rect 618 -162 675 -161
rect 761 -159 829 -158
rect 761 -161 762 -159
rect 764 -161 829 -159
rect 761 -162 829 -161
rect 885 -159 942 -158
rect 885 -161 886 -159
rect 888 -161 939 -159
rect 941 -161 942 -159
rect 885 -162 942 -161
rect 1028 -159 1096 -158
rect 1028 -161 1029 -159
rect 1031 -161 1096 -159
rect 1028 -162 1096 -161
rect 1152 -159 1209 -158
rect 1152 -161 1153 -159
rect 1155 -161 1206 -159
rect 1208 -161 1209 -159
rect 1152 -162 1209 -161
rect 1295 -159 1363 -158
rect 1295 -161 1296 -159
rect 1298 -161 1363 -159
rect 1295 -162 1363 -161
rect 1419 -159 1476 -158
rect 1419 -161 1420 -159
rect 1422 -161 1473 -159
rect 1475 -161 1476 -159
rect 1419 -162 1476 -161
rect 1562 -159 1630 -158
rect 1562 -161 1563 -159
rect 1565 -161 1630 -159
rect 1562 -162 1630 -161
rect 1686 -159 1743 -158
rect 1686 -161 1687 -159
rect 1689 -161 1740 -159
rect 1742 -161 1743 -159
rect 1686 -162 1743 -161
rect 1829 -159 1897 -158
rect 1829 -161 1830 -159
rect 1832 -161 1897 -159
rect 1829 -162 1897 -161
rect 1968 -159 2021 -158
rect 1968 -161 1969 -159
rect 1971 -161 2018 -159
rect 2020 -161 2021 -159
rect 1968 -162 2021 -161
rect 2115 -159 2183 -158
rect 2115 -161 2116 -159
rect 2118 -161 2183 -159
rect 2235 -158 2239 -157
rect 2235 -160 2236 -158
rect 2238 -160 2239 -158
rect 2235 -161 2239 -160
rect 2299 -158 2311 -157
rect 2299 -160 2300 -158
rect 2302 -160 2308 -158
rect 2310 -160 2311 -158
rect 2299 -161 2311 -160
rect 2115 -162 2183 -161
rect 2195 -162 2239 -161
rect 2195 -164 2196 -162
rect 2198 -164 2239 -162
rect 2195 -165 2239 -164
rect 80 -167 143 -166
rect 80 -169 81 -167
rect 83 -169 140 -167
rect 142 -169 143 -167
rect 80 -170 143 -169
rect 169 -167 272 -166
rect 169 -169 170 -167
rect 172 -169 268 -167
rect 270 -169 272 -167
rect 169 -170 272 -169
rect 347 -167 410 -166
rect 347 -169 348 -167
rect 350 -169 407 -167
rect 409 -169 410 -167
rect 347 -170 410 -169
rect 436 -167 539 -166
rect 436 -169 437 -167
rect 439 -169 535 -167
rect 537 -169 539 -167
rect 436 -170 539 -169
rect 614 -167 677 -166
rect 614 -169 615 -167
rect 617 -169 674 -167
rect 676 -169 677 -167
rect 614 -170 677 -169
rect 703 -167 806 -166
rect 703 -169 704 -167
rect 706 -169 802 -167
rect 804 -169 806 -167
rect 703 -170 806 -169
rect 881 -167 944 -166
rect 881 -169 882 -167
rect 884 -169 941 -167
rect 943 -169 944 -167
rect 881 -170 944 -169
rect 970 -167 1073 -166
rect 970 -169 971 -167
rect 973 -169 1069 -167
rect 1071 -169 1073 -167
rect 970 -170 1073 -169
rect 1148 -167 1211 -166
rect 1148 -169 1149 -167
rect 1151 -169 1208 -167
rect 1210 -169 1211 -167
rect 1148 -170 1211 -169
rect 1237 -167 1340 -166
rect 1237 -169 1238 -167
rect 1240 -169 1336 -167
rect 1338 -169 1340 -167
rect 1237 -170 1340 -169
rect 1415 -167 1478 -166
rect 1415 -169 1416 -167
rect 1418 -169 1475 -167
rect 1477 -169 1478 -167
rect 1415 -170 1478 -169
rect 1504 -167 1607 -166
rect 1504 -169 1505 -167
rect 1507 -169 1603 -167
rect 1605 -169 1607 -167
rect 1504 -170 1607 -169
rect 1682 -167 1745 -166
rect 1682 -169 1683 -167
rect 1685 -169 1742 -167
rect 1744 -169 1745 -167
rect 1682 -170 1745 -169
rect 1771 -167 1874 -166
rect 1771 -169 1772 -167
rect 1774 -169 1870 -167
rect 1872 -169 1874 -167
rect 1771 -170 1874 -169
rect 2057 -167 2160 -166
rect 2057 -169 2058 -167
rect 2060 -169 2156 -167
rect 2158 -169 2160 -167
rect 2057 -170 2160 -169
rect 299 -171 307 -170
rect 566 -171 574 -170
rect 833 -171 841 -170
rect 1100 -171 1108 -170
rect 1367 -171 1375 -170
rect 1634 -171 1642 -170
rect 1901 -171 1909 -170
rect 44 -172 60 -171
rect 44 -174 45 -172
rect 47 -174 57 -172
rect 59 -174 60 -172
rect 299 -173 300 -171
rect 302 -173 304 -171
rect 306 -173 307 -171
rect 299 -174 307 -173
rect 311 -172 327 -171
rect 311 -174 312 -172
rect 314 -174 324 -172
rect 326 -174 327 -172
rect 566 -173 567 -171
rect 569 -173 571 -171
rect 573 -173 574 -171
rect 566 -174 574 -173
rect 578 -172 594 -171
rect 578 -174 579 -172
rect 581 -174 591 -172
rect 593 -174 594 -172
rect 833 -173 834 -171
rect 836 -173 838 -171
rect 840 -173 841 -171
rect 833 -174 841 -173
rect 845 -172 861 -171
rect 845 -174 846 -172
rect 848 -174 858 -172
rect 860 -174 861 -172
rect 1100 -173 1101 -171
rect 1103 -173 1105 -171
rect 1107 -173 1108 -171
rect 1100 -174 1108 -173
rect 1112 -172 1128 -171
rect 1112 -174 1113 -172
rect 1115 -174 1125 -172
rect 1127 -174 1128 -172
rect 1367 -173 1368 -171
rect 1370 -173 1372 -171
rect 1374 -173 1375 -171
rect 1367 -174 1375 -173
rect 1379 -172 1395 -171
rect 1379 -174 1380 -172
rect 1382 -174 1392 -172
rect 1394 -174 1395 -172
rect 1634 -173 1635 -171
rect 1637 -173 1639 -171
rect 1641 -173 1642 -171
rect 1634 -174 1642 -173
rect 1646 -172 1662 -171
rect 1646 -174 1647 -172
rect 1649 -174 1659 -172
rect 1661 -174 1662 -172
rect 1901 -173 1902 -171
rect 1904 -173 1906 -171
rect 1908 -173 1909 -171
rect 1901 -174 1909 -173
rect 2187 -171 2195 -170
rect 2187 -173 2188 -171
rect 2190 -173 2192 -171
rect 2194 -173 2195 -171
rect 2187 -174 2195 -173
rect 44 -175 60 -174
rect 88 -175 214 -174
rect 311 -175 327 -174
rect 355 -175 481 -174
rect 578 -175 594 -174
rect 622 -175 748 -174
rect 845 -175 861 -174
rect 889 -175 1015 -174
rect 1112 -175 1128 -174
rect 1156 -175 1282 -174
rect 1379 -175 1395 -174
rect 1423 -175 1549 -174
rect 1646 -175 1662 -174
rect 1690 -175 1816 -174
rect 1976 -175 2102 -174
rect 88 -177 89 -175
rect 91 -177 211 -175
rect 213 -177 214 -175
rect 88 -178 214 -177
rect 355 -177 356 -175
rect 358 -177 478 -175
rect 480 -177 481 -175
rect 355 -178 481 -177
rect 622 -177 623 -175
rect 625 -177 745 -175
rect 747 -177 748 -175
rect 622 -178 748 -177
rect 889 -177 890 -175
rect 892 -177 1012 -175
rect 1014 -177 1015 -175
rect 889 -178 1015 -177
rect 1156 -177 1157 -175
rect 1159 -177 1279 -175
rect 1281 -177 1282 -175
rect 1156 -178 1282 -177
rect 1423 -177 1424 -175
rect 1426 -177 1546 -175
rect 1548 -177 1549 -175
rect 1423 -178 1549 -177
rect 1690 -177 1691 -175
rect 1693 -177 1813 -175
rect 1815 -177 1816 -175
rect 1690 -178 1816 -177
rect 1840 -176 1864 -175
rect 1840 -178 1841 -176
rect 1843 -178 1861 -176
rect 1863 -178 1864 -176
rect 1840 -179 1864 -178
rect 1924 -176 1932 -175
rect 1924 -178 1925 -176
rect 1927 -178 1929 -176
rect 1931 -178 1932 -176
rect 1976 -177 1977 -175
rect 1979 -177 2099 -175
rect 2101 -177 2102 -175
rect 1976 -178 2102 -177
rect 2209 -175 2213 -174
rect 2209 -177 2210 -175
rect 2212 -177 2213 -175
rect 2209 -178 2213 -177
rect 1924 -179 1932 -178
rect 2146 -179 2213 -178
rect 2146 -181 2147 -179
rect 2149 -181 2213 -179
rect 2146 -182 2213 -181
rect 2275 -175 2279 -174
rect 2275 -177 2276 -175
rect 2278 -177 2279 -175
rect 260 -184 339 -183
rect 260 -186 261 -184
rect 263 -186 336 -184
rect 338 -186 339 -184
rect 260 -187 339 -186
rect 527 -184 606 -183
rect 527 -186 528 -184
rect 530 -186 603 -184
rect 605 -186 606 -184
rect 527 -187 606 -186
rect 794 -184 873 -183
rect 794 -186 795 -184
rect 797 -186 870 -184
rect 872 -186 873 -184
rect 794 -187 873 -186
rect 1061 -184 1140 -183
rect 1061 -186 1062 -184
rect 1064 -186 1137 -184
rect 1139 -186 1140 -184
rect 1061 -187 1140 -186
rect 1328 -184 1407 -183
rect 1328 -186 1329 -184
rect 1331 -186 1404 -184
rect 1406 -186 1407 -184
rect 1328 -187 1407 -186
rect 1595 -184 1674 -183
rect 1595 -186 1596 -184
rect 1598 -186 1671 -184
rect 1673 -186 1674 -184
rect 1595 -187 1674 -186
rect 2275 -199 2279 -177
rect 2323 -193 2331 -192
rect 2323 -195 2324 -193
rect 2326 -195 2328 -193
rect 2330 -195 2331 -193
rect 2323 -196 2331 -195
rect 2275 -201 2276 -199
rect 2278 -201 2279 -199
rect 128 -202 136 -201
rect 128 -204 129 -202
rect 131 -204 133 -202
rect 135 -204 136 -202
rect 128 -205 136 -204
rect 395 -202 403 -201
rect 395 -204 400 -202
rect 402 -204 403 -202
rect 395 -205 403 -204
rect 662 -202 670 -201
rect 662 -204 667 -202
rect 669 -204 670 -202
rect 662 -205 670 -204
rect 929 -202 937 -201
rect 929 -204 934 -202
rect 936 -204 937 -202
rect 929 -205 937 -204
rect 1196 -202 1204 -201
rect 1196 -204 1201 -202
rect 1203 -204 1204 -202
rect 1196 -205 1204 -204
rect 1463 -202 1471 -201
rect 1463 -204 1468 -202
rect 1470 -204 1471 -202
rect 1463 -205 1471 -204
rect 1730 -202 1738 -201
rect 1730 -204 1735 -202
rect 1737 -204 1738 -202
rect 1730 -205 1738 -204
rect 260 -214 355 -213
rect 260 -216 261 -214
rect 263 -216 352 -214
rect 354 -216 355 -214
rect 260 -217 355 -216
rect 527 -214 622 -213
rect 527 -216 528 -214
rect 530 -216 619 -214
rect 621 -216 622 -214
rect 527 -217 622 -216
rect 794 -214 889 -213
rect 794 -216 795 -214
rect 797 -216 886 -214
rect 888 -216 889 -214
rect 794 -217 889 -216
rect 1061 -214 1156 -213
rect 1061 -216 1062 -214
rect 1064 -216 1153 -214
rect 1155 -216 1156 -214
rect 1061 -217 1156 -216
rect 1328 -214 1423 -213
rect 1328 -216 1329 -214
rect 1331 -216 1420 -214
rect 1422 -216 1423 -214
rect 1328 -217 1423 -216
rect 1595 -214 1690 -213
rect 1595 -216 1596 -214
rect 1598 -216 1687 -214
rect 1689 -216 1690 -214
rect 1595 -217 1690 -216
rect 1862 -214 1892 -213
rect 1862 -216 1863 -214
rect 1865 -216 1889 -214
rect 1891 -216 1892 -214
rect 1862 -217 1892 -216
rect 2148 -214 2213 -213
rect 2148 -216 2149 -214
rect 2151 -216 2213 -214
rect 2148 -217 2213 -216
rect 1924 -222 1932 -221
rect 88 -223 214 -222
rect 88 -225 89 -223
rect 91 -225 211 -223
rect 213 -225 214 -223
rect 355 -223 481 -222
rect 88 -226 214 -225
rect 218 -225 271 -224
rect 218 -227 268 -225
rect 270 -227 271 -225
rect 355 -225 356 -223
rect 358 -225 478 -223
rect 480 -225 481 -223
rect 622 -223 748 -222
rect 355 -226 481 -225
rect 485 -225 538 -224
rect 218 -228 271 -227
rect 485 -227 535 -225
rect 537 -227 538 -225
rect 622 -225 623 -223
rect 625 -225 745 -223
rect 747 -225 748 -223
rect 889 -223 1015 -222
rect 622 -226 748 -225
rect 752 -225 805 -224
rect 485 -228 538 -227
rect 752 -227 802 -225
rect 804 -227 805 -225
rect 889 -225 890 -223
rect 892 -225 1012 -223
rect 1014 -225 1015 -223
rect 1156 -223 1282 -222
rect 889 -226 1015 -225
rect 1019 -225 1072 -224
rect 752 -228 805 -227
rect 1019 -227 1069 -225
rect 1071 -227 1072 -225
rect 1156 -225 1157 -223
rect 1159 -225 1279 -223
rect 1281 -225 1282 -223
rect 1423 -223 1549 -222
rect 1156 -226 1282 -225
rect 1286 -225 1339 -224
rect 1019 -228 1072 -227
rect 1286 -227 1336 -225
rect 1338 -227 1339 -225
rect 1423 -225 1424 -223
rect 1426 -225 1546 -223
rect 1548 -225 1549 -223
rect 1690 -223 1816 -222
rect 1423 -226 1549 -225
rect 1553 -225 1606 -224
rect 1286 -228 1339 -227
rect 1553 -227 1603 -225
rect 1605 -227 1606 -225
rect 1690 -225 1691 -223
rect 1693 -225 1813 -223
rect 1815 -225 1816 -223
rect 1924 -224 1925 -222
rect 1927 -224 1929 -222
rect 1931 -224 1932 -222
rect 1690 -226 1816 -225
rect 1820 -225 1873 -224
rect 1924 -225 1932 -224
rect 1976 -223 2102 -222
rect 1976 -225 1977 -223
rect 1979 -225 2099 -223
rect 2101 -225 2102 -223
rect 2209 -223 2213 -217
rect 1553 -228 1606 -227
rect 1820 -227 1870 -225
rect 1872 -227 1873 -225
rect 1976 -226 2102 -225
rect 2106 -225 2159 -224
rect 1820 -228 1873 -227
rect 2106 -227 2156 -225
rect 2158 -227 2159 -225
rect 2209 -225 2210 -223
rect 2212 -225 2213 -223
rect 2209 -226 2213 -225
rect 2275 -223 2279 -201
rect 2275 -225 2276 -223
rect 2278 -225 2279 -223
rect 2275 -226 2279 -225
rect 2106 -228 2159 -227
rect 2187 -228 2203 -227
rect 218 -230 222 -228
rect 485 -230 489 -228
rect 752 -230 756 -228
rect 1019 -230 1023 -228
rect 1286 -230 1290 -228
rect 1553 -230 1557 -228
rect 1820 -230 1824 -228
rect 2106 -230 2110 -228
rect 36 -231 44 -230
rect 36 -233 37 -231
rect 39 -233 41 -231
rect 43 -233 44 -231
rect 36 -234 44 -233
rect 80 -231 142 -230
rect 80 -233 81 -231
rect 83 -233 139 -231
rect 141 -233 142 -231
rect 80 -234 142 -233
rect 169 -231 222 -230
rect 169 -233 170 -231
rect 172 -233 222 -231
rect 169 -234 222 -233
rect 347 -231 409 -230
rect 347 -233 348 -231
rect 350 -233 406 -231
rect 408 -233 409 -231
rect 347 -234 409 -233
rect 436 -231 489 -230
rect 436 -233 437 -231
rect 439 -233 489 -231
rect 436 -234 489 -233
rect 614 -231 676 -230
rect 614 -233 615 -231
rect 617 -233 673 -231
rect 675 -233 676 -231
rect 614 -234 676 -233
rect 703 -231 756 -230
rect 703 -233 704 -231
rect 706 -233 756 -231
rect 703 -234 756 -233
rect 881 -231 943 -230
rect 881 -233 882 -231
rect 884 -233 940 -231
rect 942 -233 943 -231
rect 881 -234 943 -233
rect 970 -231 1023 -230
rect 970 -233 971 -231
rect 973 -233 1023 -231
rect 970 -234 1023 -233
rect 1148 -231 1210 -230
rect 1148 -233 1149 -231
rect 1151 -233 1207 -231
rect 1209 -233 1210 -231
rect 1148 -234 1210 -233
rect 1237 -231 1290 -230
rect 1237 -233 1238 -231
rect 1240 -233 1290 -231
rect 1237 -234 1290 -233
rect 1415 -231 1477 -230
rect 1415 -233 1416 -231
rect 1418 -233 1474 -231
rect 1476 -233 1477 -231
rect 1415 -234 1477 -233
rect 1504 -231 1557 -230
rect 1504 -233 1505 -231
rect 1507 -233 1557 -231
rect 1504 -234 1557 -233
rect 1682 -231 1744 -230
rect 1682 -233 1683 -231
rect 1685 -233 1741 -231
rect 1743 -233 1744 -231
rect 1682 -234 1744 -233
rect 1771 -231 1824 -230
rect 1771 -233 1772 -231
rect 1774 -233 1824 -231
rect 1771 -234 1824 -233
rect 2057 -231 2110 -230
rect 2187 -230 2188 -228
rect 2190 -230 2200 -228
rect 2202 -230 2203 -228
rect 2187 -231 2203 -230
rect 2057 -233 2058 -231
rect 2060 -233 2110 -231
rect 2057 -234 2110 -233
rect 227 -236 307 -235
rect 227 -238 228 -236
rect 230 -238 304 -236
rect 306 -238 307 -236
rect 494 -236 574 -235
rect 494 -238 495 -236
rect 497 -238 571 -236
rect 573 -238 574 -236
rect 761 -236 841 -235
rect 761 -238 762 -236
rect 764 -238 838 -236
rect 840 -238 841 -236
rect 1028 -236 1108 -235
rect 1028 -238 1029 -236
rect 1031 -238 1105 -236
rect 1107 -238 1108 -236
rect 1295 -236 1375 -235
rect 1295 -238 1296 -236
rect 1298 -238 1372 -236
rect 1374 -238 1375 -236
rect 1562 -236 1642 -235
rect 1562 -238 1563 -236
rect 1565 -238 1639 -236
rect 1641 -238 1642 -236
rect 1829 -236 1909 -235
rect 1829 -238 1830 -236
rect 1832 -238 1906 -236
rect 1908 -238 1909 -236
rect 2115 -236 2195 -235
rect 2115 -238 2116 -236
rect 2118 -238 2192 -236
rect 2194 -238 2195 -236
rect 128 -239 136 -238
rect 227 -239 307 -238
rect 395 -239 403 -238
rect 494 -239 574 -238
rect 662 -239 670 -238
rect 761 -239 841 -238
rect 929 -239 937 -238
rect 1028 -239 1108 -238
rect 1196 -239 1204 -238
rect 1295 -239 1375 -238
rect 1463 -239 1471 -238
rect 1562 -239 1642 -238
rect 1730 -239 1738 -238
rect 1829 -239 1909 -238
rect 1968 -239 2021 -238
rect 2115 -239 2195 -238
rect 2299 -238 2323 -237
rect 128 -241 129 -239
rect 131 -241 133 -239
rect 135 -241 136 -239
rect 128 -242 136 -241
rect 395 -241 396 -239
rect 398 -241 400 -239
rect 402 -241 403 -239
rect 395 -242 403 -241
rect 662 -241 663 -239
rect 665 -241 667 -239
rect 669 -241 670 -239
rect 662 -242 670 -241
rect 929 -241 930 -239
rect 932 -241 934 -239
rect 936 -241 937 -239
rect 929 -242 937 -241
rect 1196 -241 1197 -239
rect 1199 -241 1201 -239
rect 1203 -241 1204 -239
rect 1196 -242 1204 -241
rect 1463 -241 1464 -239
rect 1466 -241 1468 -239
rect 1470 -241 1471 -239
rect 1463 -242 1471 -241
rect 1730 -241 1731 -239
rect 1733 -241 1735 -239
rect 1737 -241 1738 -239
rect 1730 -242 1738 -241
rect 1968 -241 1969 -239
rect 1971 -241 2018 -239
rect 2020 -241 2021 -239
rect 1968 -242 2021 -241
rect 2235 -240 2247 -239
rect 2235 -242 2236 -240
rect 2238 -242 2244 -240
rect 2246 -242 2247 -240
rect 2299 -240 2300 -238
rect 2302 -240 2320 -238
rect 2322 -240 2323 -238
rect 2299 -241 2323 -240
rect 2 -243 12 -242
rect 2235 -243 2247 -242
rect 2 -245 3 -243
rect 5 -245 9 -243
rect 11 -245 12 -243
rect 2 -246 12 -245
rect 44 -244 52 -243
rect 44 -246 45 -244
rect 47 -246 49 -244
rect 51 -246 52 -244
rect 44 -247 52 -246
rect 179 -244 271 -243
rect 179 -246 180 -244
rect 182 -246 268 -244
rect 270 -246 271 -244
rect 179 -247 271 -246
rect 311 -244 319 -243
rect 311 -246 312 -244
rect 314 -246 316 -244
rect 318 -246 319 -244
rect 311 -247 319 -246
rect 446 -244 538 -243
rect 446 -246 447 -244
rect 449 -246 535 -244
rect 537 -246 538 -244
rect 446 -247 538 -246
rect 578 -244 586 -243
rect 578 -246 579 -244
rect 581 -246 583 -244
rect 585 -246 586 -244
rect 578 -247 586 -246
rect 713 -244 805 -243
rect 713 -246 714 -244
rect 716 -246 802 -244
rect 804 -246 805 -244
rect 713 -247 805 -246
rect 845 -244 853 -243
rect 845 -246 846 -244
rect 848 -246 850 -244
rect 852 -246 853 -244
rect 845 -247 853 -246
rect 980 -244 1072 -243
rect 980 -246 981 -244
rect 983 -246 1069 -244
rect 1071 -246 1072 -244
rect 980 -247 1072 -246
rect 1112 -244 1120 -243
rect 1112 -246 1113 -244
rect 1115 -246 1117 -244
rect 1119 -246 1120 -244
rect 1112 -247 1120 -246
rect 1247 -244 1339 -243
rect 1247 -246 1248 -244
rect 1250 -246 1336 -244
rect 1338 -246 1339 -244
rect 1247 -247 1339 -246
rect 1379 -244 1387 -243
rect 1379 -246 1380 -244
rect 1382 -246 1384 -244
rect 1386 -246 1387 -244
rect 1379 -247 1387 -246
rect 1514 -244 1606 -243
rect 1514 -246 1515 -244
rect 1517 -246 1603 -244
rect 1605 -246 1606 -244
rect 1514 -247 1606 -246
rect 1646 -244 1654 -243
rect 1646 -246 1647 -244
rect 1649 -246 1651 -244
rect 1653 -246 1654 -244
rect 1646 -247 1654 -246
rect 1781 -244 1873 -243
rect 1781 -246 1782 -244
rect 1784 -246 1870 -244
rect 1872 -246 1873 -244
rect 1781 -247 1873 -246
rect 2067 -244 2159 -243
rect 2067 -246 2068 -244
rect 2070 -246 2156 -244
rect 2158 -246 2159 -244
rect 2067 -247 2159 -246
rect 299 -256 400 -255
rect 299 -258 300 -256
rect 302 -258 396 -256
rect 398 -258 400 -256
rect 299 -259 400 -258
rect 566 -256 667 -255
rect 566 -258 567 -256
rect 569 -258 663 -256
rect 665 -258 667 -256
rect 566 -259 667 -258
rect 833 -256 934 -255
rect 833 -258 834 -256
rect 836 -258 930 -256
rect 932 -258 934 -256
rect 833 -259 934 -258
rect 1100 -256 1201 -255
rect 1100 -258 1101 -256
rect 1103 -258 1197 -256
rect 1199 -258 1201 -256
rect 1100 -259 1201 -258
rect 1367 -256 1468 -255
rect 1367 -258 1368 -256
rect 1370 -258 1464 -256
rect 1466 -258 1468 -256
rect 1367 -259 1468 -258
rect 1634 -256 1735 -255
rect 1634 -258 1635 -256
rect 1637 -258 1731 -256
rect 1733 -258 1735 -256
rect 1634 -259 1735 -258
rect 1896 -256 1905 -255
rect 1896 -258 1897 -256
rect 1899 -258 1902 -256
rect 1904 -258 1905 -256
rect 1896 -259 1905 -258
rect 2327 -265 2331 -264
rect 2327 -267 2328 -265
rect 2330 -267 2331 -265
rect 2327 -269 2331 -267
rect 2327 -271 2328 -269
rect 2330 -271 2331 -269
rect 2327 -272 2331 -271
<< alu3 >>
rect 1769 300 2196 304
rect 262 286 266 287
rect 262 284 263 286
rect 265 284 266 286
rect 2 276 6 277
rect 2 274 3 276
rect 5 274 6 276
rect 262 274 266 284
rect 529 278 533 279
rect 529 276 530 278
rect 532 276 533 278
rect 2 205 6 274
rect 212 273 216 274
rect 212 271 213 273
rect 215 271 216 273
rect 262 272 263 274
rect 265 272 266 274
rect 262 271 266 272
rect 351 273 355 274
rect 351 271 352 273
rect 354 271 355 273
rect 2 203 3 205
rect 5 203 6 205
rect 2 132 6 203
rect 2 130 3 132
rect 5 130 6 132
rect 2 61 6 130
rect 2 59 3 61
rect 5 59 6 61
rect 2 -12 6 59
rect 2 -14 3 -12
rect 5 -14 6 -12
rect 2 -83 6 -14
rect 2 -85 3 -83
rect 5 -85 6 -83
rect 2 -156 6 -85
rect 2 -158 3 -156
rect 5 -158 6 -156
rect 2 -243 6 -158
rect 44 259 48 260
rect 44 257 45 259
rect 47 257 48 259
rect 44 185 48 257
rect 212 236 216 271
rect 212 234 213 236
rect 215 234 216 236
rect 212 233 216 234
rect 303 261 307 262
rect 303 259 304 261
rect 306 259 307 261
rect 303 196 307 259
rect 303 194 304 196
rect 306 194 307 196
rect 303 193 307 194
rect 311 259 315 260
rect 311 257 312 259
rect 314 257 315 259
rect 44 183 45 185
rect 47 183 48 185
rect 44 116 48 183
rect 311 185 315 257
rect 351 218 355 271
rect 479 273 483 274
rect 479 271 480 273
rect 482 271 483 273
rect 479 236 483 271
rect 529 273 533 276
rect 529 271 530 273
rect 532 271 533 273
rect 529 270 533 271
rect 618 273 622 274
rect 618 271 619 273
rect 621 271 622 273
rect 479 234 480 236
rect 482 234 483 236
rect 479 233 483 234
rect 570 261 574 262
rect 570 259 571 261
rect 573 259 574 261
rect 351 216 352 218
rect 354 216 355 218
rect 351 215 355 216
rect 570 196 574 259
rect 570 194 571 196
rect 573 194 574 196
rect 311 183 312 185
rect 314 183 315 185
rect 44 114 45 116
rect 47 114 48 116
rect 44 41 48 114
rect 303 117 307 118
rect 303 115 304 117
rect 306 115 307 117
rect 303 52 307 115
rect 303 50 304 52
rect 306 50 307 52
rect 303 49 307 50
rect 311 116 315 183
rect 311 114 312 116
rect 314 114 315 116
rect 44 39 45 41
rect 47 39 48 41
rect 44 -29 48 39
rect 311 41 315 114
rect 335 193 339 194
rect 570 193 574 194
rect 578 259 582 260
rect 578 257 579 259
rect 581 257 582 259
rect 335 191 336 193
rect 338 191 339 193
rect 335 104 339 191
rect 578 185 582 257
rect 618 218 622 271
rect 746 273 750 274
rect 746 271 747 273
rect 749 271 750 273
rect 885 273 889 274
rect 885 271 886 273
rect 888 271 889 273
rect 746 236 750 271
rect 796 270 800 271
rect 796 268 797 270
rect 799 268 800 270
rect 796 257 800 268
rect 796 255 797 257
rect 799 255 800 257
rect 796 254 800 255
rect 837 261 841 262
rect 837 259 838 261
rect 840 259 841 261
rect 746 234 747 236
rect 749 234 750 236
rect 746 233 750 234
rect 618 216 619 218
rect 621 216 622 218
rect 618 215 622 216
rect 837 196 841 259
rect 837 194 838 196
rect 840 194 841 196
rect 578 183 579 185
rect 581 183 582 185
rect 335 102 336 104
rect 338 102 339 104
rect 335 101 339 102
rect 351 129 355 130
rect 351 127 352 129
rect 354 127 355 129
rect 351 74 355 127
rect 351 72 352 74
rect 354 72 355 74
rect 351 71 355 72
rect 570 117 574 118
rect 570 115 571 117
rect 573 115 574 117
rect 570 52 574 115
rect 570 50 571 52
rect 573 50 574 52
rect 311 39 312 41
rect 314 39 315 41
rect 44 -31 45 -29
rect 47 -31 48 -29
rect 44 -103 48 -31
rect 303 -27 307 -26
rect 303 -29 304 -27
rect 306 -29 307 -27
rect 303 -92 307 -29
rect 303 -94 304 -92
rect 306 -94 307 -92
rect 303 -95 307 -94
rect 311 -29 315 39
rect 311 -31 312 -29
rect 314 -31 315 -29
rect 44 -105 45 -103
rect 47 -105 48 -103
rect 44 -172 48 -105
rect 311 -103 315 -31
rect 335 49 339 50
rect 570 49 574 50
rect 578 116 582 183
rect 578 114 579 116
rect 581 114 582 116
rect 335 47 336 49
rect 338 47 339 49
rect 335 -40 339 47
rect 578 41 582 114
rect 602 193 606 194
rect 837 193 841 194
rect 845 259 849 260
rect 845 257 846 259
rect 848 257 849 259
rect 602 191 603 193
rect 605 191 606 193
rect 602 104 606 191
rect 845 185 849 257
rect 885 218 889 271
rect 1013 273 1017 274
rect 1013 271 1014 273
rect 1016 271 1017 273
rect 1013 236 1017 271
rect 1152 273 1156 274
rect 1152 271 1153 273
rect 1155 271 1156 273
rect 1063 262 1067 263
rect 1063 260 1064 262
rect 1066 260 1067 262
rect 1063 257 1067 260
rect 1063 255 1064 257
rect 1066 255 1067 257
rect 1063 254 1067 255
rect 1104 261 1108 262
rect 1104 259 1105 261
rect 1107 259 1108 261
rect 1013 234 1014 236
rect 1016 234 1017 236
rect 1013 233 1017 234
rect 885 216 886 218
rect 888 216 889 218
rect 885 215 889 216
rect 1104 196 1108 259
rect 1104 194 1105 196
rect 1107 194 1108 196
rect 845 183 846 185
rect 848 183 849 185
rect 602 102 603 104
rect 605 102 606 104
rect 602 101 606 102
rect 618 129 622 130
rect 618 127 619 129
rect 621 127 622 129
rect 618 74 622 127
rect 618 72 619 74
rect 621 72 622 74
rect 618 71 622 72
rect 837 117 841 118
rect 837 115 838 117
rect 840 115 841 117
rect 837 52 841 115
rect 837 50 838 52
rect 840 50 841 52
rect 578 39 579 41
rect 581 39 582 41
rect 335 -42 336 -40
rect 338 -42 339 -40
rect 335 -43 339 -42
rect 351 -15 355 -14
rect 351 -17 352 -15
rect 354 -17 355 -15
rect 351 -70 355 -17
rect 351 -72 352 -70
rect 354 -72 355 -70
rect 351 -73 355 -72
rect 570 -27 574 -26
rect 570 -29 571 -27
rect 573 -29 574 -27
rect 570 -92 574 -29
rect 570 -94 571 -92
rect 573 -94 574 -92
rect 311 -105 312 -103
rect 314 -105 315 -103
rect 44 -174 45 -172
rect 47 -174 48 -172
rect 36 -231 40 -230
rect 36 -233 37 -231
rect 39 -233 40 -231
rect 36 -236 40 -233
rect 36 -238 37 -236
rect 39 -238 40 -236
rect 36 -239 40 -238
rect 2 -245 3 -243
rect 5 -245 6 -243
rect 2 -249 6 -245
rect 44 -244 48 -174
rect 303 -171 307 -170
rect 303 -173 304 -171
rect 306 -173 307 -171
rect 128 -202 132 -201
rect 128 -204 129 -202
rect 131 -204 132 -202
rect 128 -239 132 -204
rect 303 -236 307 -173
rect 303 -238 304 -236
rect 306 -238 307 -236
rect 303 -239 307 -238
rect 311 -172 315 -105
rect 311 -174 312 -172
rect 314 -174 315 -172
rect 128 -241 129 -239
rect 131 -241 132 -239
rect 128 -242 132 -241
rect 44 -246 45 -244
rect 47 -246 48 -244
rect 44 -247 48 -246
rect 311 -244 315 -174
rect 335 -95 339 -94
rect 570 -95 574 -94
rect 578 -29 582 39
rect 578 -31 579 -29
rect 581 -31 582 -29
rect 335 -97 336 -95
rect 338 -97 339 -95
rect 335 -184 339 -97
rect 578 -103 582 -31
rect 602 49 606 50
rect 837 49 841 50
rect 845 116 849 183
rect 845 114 846 116
rect 848 114 849 116
rect 602 47 603 49
rect 605 47 606 49
rect 602 -40 606 47
rect 845 41 849 114
rect 869 193 873 194
rect 1104 193 1108 194
rect 1112 259 1116 260
rect 1112 257 1113 259
rect 1115 257 1116 259
rect 869 191 870 193
rect 872 191 873 193
rect 869 104 873 191
rect 1112 185 1116 257
rect 1152 218 1156 271
rect 1280 273 1284 274
rect 1280 271 1281 273
rect 1283 271 1284 273
rect 1280 236 1284 271
rect 1419 273 1423 274
rect 1419 271 1420 273
rect 1422 271 1423 273
rect 1371 261 1375 262
rect 1371 259 1372 261
rect 1374 259 1375 261
rect 1330 254 1334 255
rect 1330 252 1331 254
rect 1333 252 1334 254
rect 1330 248 1334 252
rect 1330 246 1331 248
rect 1333 246 1334 248
rect 1330 245 1334 246
rect 1280 234 1281 236
rect 1283 234 1284 236
rect 1280 233 1284 234
rect 1152 216 1153 218
rect 1155 216 1156 218
rect 1152 215 1156 216
rect 1371 196 1375 259
rect 1371 194 1372 196
rect 1374 194 1375 196
rect 1112 183 1113 185
rect 1115 183 1116 185
rect 869 102 870 104
rect 872 102 873 104
rect 869 101 873 102
rect 885 129 889 130
rect 885 127 886 129
rect 888 127 889 129
rect 885 74 889 127
rect 885 72 886 74
rect 888 72 889 74
rect 885 71 889 72
rect 1104 117 1108 118
rect 1104 115 1105 117
rect 1107 115 1108 117
rect 1104 52 1108 115
rect 1104 50 1105 52
rect 1107 50 1108 52
rect 845 39 846 41
rect 848 39 849 41
rect 602 -42 603 -40
rect 605 -42 606 -40
rect 602 -43 606 -42
rect 618 -15 622 -14
rect 618 -17 619 -15
rect 621 -17 622 -15
rect 618 -70 622 -17
rect 618 -72 619 -70
rect 621 -72 622 -70
rect 618 -73 622 -72
rect 837 -27 841 -26
rect 837 -29 838 -27
rect 840 -29 841 -27
rect 837 -92 841 -29
rect 837 -94 838 -92
rect 840 -94 841 -92
rect 578 -105 579 -103
rect 581 -105 582 -103
rect 335 -186 336 -184
rect 338 -186 339 -184
rect 335 -187 339 -186
rect 351 -159 355 -158
rect 351 -161 352 -159
rect 354 -161 355 -159
rect 351 -214 355 -161
rect 351 -216 352 -214
rect 354 -216 355 -214
rect 351 -217 355 -216
rect 570 -171 574 -170
rect 570 -173 571 -171
rect 573 -173 574 -171
rect 570 -236 574 -173
rect 570 -238 571 -236
rect 573 -238 574 -236
rect 311 -246 312 -244
rect 314 -246 315 -244
rect 311 -247 315 -246
rect 395 -239 399 -238
rect 570 -239 574 -238
rect 578 -172 582 -105
rect 578 -174 579 -172
rect 581 -174 582 -172
rect 395 -241 396 -239
rect 398 -241 399 -239
rect 395 -256 399 -241
rect 578 -244 582 -174
rect 602 -95 606 -94
rect 837 -95 841 -94
rect 845 -29 849 39
rect 845 -31 846 -29
rect 848 -31 849 -29
rect 602 -97 603 -95
rect 605 -97 606 -95
rect 602 -184 606 -97
rect 845 -103 849 -31
rect 869 49 873 50
rect 1104 49 1108 50
rect 1112 116 1116 183
rect 1112 114 1113 116
rect 1115 114 1116 116
rect 869 47 870 49
rect 872 47 873 49
rect 869 -40 873 47
rect 1112 41 1116 114
rect 1136 193 1140 194
rect 1371 193 1375 194
rect 1379 259 1383 260
rect 1379 257 1380 259
rect 1382 257 1383 259
rect 1136 191 1137 193
rect 1139 191 1140 193
rect 1136 104 1140 191
rect 1379 185 1383 257
rect 1419 218 1423 271
rect 1547 273 1551 274
rect 1547 271 1548 273
rect 1550 271 1551 273
rect 1547 236 1551 271
rect 1686 273 1690 274
rect 1686 271 1687 273
rect 1689 271 1690 273
rect 1638 261 1642 262
rect 1638 259 1639 261
rect 1641 259 1642 261
rect 1597 250 1601 251
rect 1597 248 1598 250
rect 1600 248 1601 250
rect 1597 246 1601 248
rect 1597 244 1598 246
rect 1600 244 1601 246
rect 1597 243 1601 244
rect 1547 234 1548 236
rect 1550 234 1551 236
rect 1547 233 1551 234
rect 1419 216 1420 218
rect 1422 216 1423 218
rect 1419 215 1423 216
rect 1638 196 1642 259
rect 1638 194 1639 196
rect 1641 194 1642 196
rect 1379 183 1380 185
rect 1382 183 1383 185
rect 1136 102 1137 104
rect 1139 102 1140 104
rect 1136 101 1140 102
rect 1152 129 1156 130
rect 1152 127 1153 129
rect 1155 127 1156 129
rect 1152 74 1156 127
rect 1152 72 1153 74
rect 1155 72 1156 74
rect 1152 71 1156 72
rect 1371 117 1375 118
rect 1371 115 1372 117
rect 1374 115 1375 117
rect 1371 52 1375 115
rect 1371 50 1372 52
rect 1374 50 1375 52
rect 1112 39 1113 41
rect 1115 39 1116 41
rect 869 -42 870 -40
rect 872 -42 873 -40
rect 869 -43 873 -42
rect 885 -15 889 -14
rect 885 -17 886 -15
rect 888 -17 889 -15
rect 885 -70 889 -17
rect 885 -72 886 -70
rect 888 -72 889 -70
rect 885 -73 889 -72
rect 1104 -27 1108 -26
rect 1104 -29 1105 -27
rect 1107 -29 1108 -27
rect 1104 -92 1108 -29
rect 1104 -94 1105 -92
rect 1107 -94 1108 -92
rect 845 -105 846 -103
rect 848 -105 849 -103
rect 602 -186 603 -184
rect 605 -186 606 -184
rect 602 -187 606 -186
rect 618 -159 622 -158
rect 618 -161 619 -159
rect 621 -161 622 -159
rect 618 -214 622 -161
rect 618 -216 619 -214
rect 621 -216 622 -214
rect 618 -217 622 -216
rect 837 -171 841 -170
rect 837 -173 838 -171
rect 840 -173 841 -171
rect 837 -236 841 -173
rect 837 -238 838 -236
rect 840 -238 841 -236
rect 578 -246 579 -244
rect 581 -246 582 -244
rect 578 -247 582 -246
rect 662 -239 666 -238
rect 837 -239 841 -238
rect 845 -172 849 -105
rect 845 -174 846 -172
rect 848 -174 849 -172
rect 662 -241 663 -239
rect 665 -241 666 -239
rect 395 -258 396 -256
rect 398 -258 399 -256
rect 395 -259 399 -258
rect 662 -256 666 -241
rect 845 -244 849 -174
rect 869 -95 873 -94
rect 1104 -95 1108 -94
rect 1112 -29 1116 39
rect 1112 -31 1113 -29
rect 1115 -31 1116 -29
rect 869 -97 870 -95
rect 872 -97 873 -95
rect 869 -184 873 -97
rect 1112 -103 1116 -31
rect 1136 49 1140 50
rect 1371 49 1375 50
rect 1379 116 1383 183
rect 1379 114 1380 116
rect 1382 114 1383 116
rect 1136 47 1137 49
rect 1139 47 1140 49
rect 1136 -40 1140 47
rect 1379 41 1383 114
rect 1403 193 1407 194
rect 1638 193 1642 194
rect 1646 259 1650 260
rect 1646 257 1647 259
rect 1649 257 1650 259
rect 1403 191 1404 193
rect 1406 191 1407 193
rect 1403 104 1407 191
rect 1646 185 1650 257
rect 1686 218 1690 271
rect 1686 216 1687 218
rect 1689 216 1690 218
rect 1686 215 1690 216
rect 1646 183 1647 185
rect 1649 183 1650 185
rect 1403 102 1404 104
rect 1406 102 1407 104
rect 1403 101 1407 102
rect 1419 129 1423 130
rect 1419 127 1420 129
rect 1422 127 1423 129
rect 1419 74 1423 127
rect 1419 72 1420 74
rect 1422 72 1423 74
rect 1419 71 1423 72
rect 1638 117 1642 118
rect 1638 115 1639 117
rect 1641 115 1642 117
rect 1638 52 1642 115
rect 1638 50 1639 52
rect 1641 50 1642 52
rect 1379 39 1380 41
rect 1382 39 1383 41
rect 1136 -42 1137 -40
rect 1139 -42 1140 -40
rect 1136 -43 1140 -42
rect 1152 -15 1156 -14
rect 1152 -17 1153 -15
rect 1155 -17 1156 -15
rect 1152 -70 1156 -17
rect 1152 -72 1153 -70
rect 1155 -72 1156 -70
rect 1152 -73 1156 -72
rect 1371 -27 1375 -26
rect 1371 -29 1372 -27
rect 1374 -29 1375 -27
rect 1371 -92 1375 -29
rect 1371 -94 1372 -92
rect 1374 -94 1375 -92
rect 1112 -105 1113 -103
rect 1115 -105 1116 -103
rect 869 -186 870 -184
rect 872 -186 873 -184
rect 869 -187 873 -186
rect 885 -159 889 -158
rect 885 -161 886 -159
rect 888 -161 889 -159
rect 885 -214 889 -161
rect 885 -216 886 -214
rect 888 -216 889 -214
rect 885 -217 889 -216
rect 1104 -171 1108 -170
rect 1104 -173 1105 -171
rect 1107 -173 1108 -171
rect 1104 -236 1108 -173
rect 1104 -238 1105 -236
rect 1107 -238 1108 -236
rect 845 -246 846 -244
rect 848 -246 849 -244
rect 845 -247 849 -246
rect 929 -239 933 -238
rect 1104 -239 1108 -238
rect 1112 -172 1116 -105
rect 1112 -174 1113 -172
rect 1115 -174 1116 -172
rect 929 -241 930 -239
rect 932 -241 933 -239
rect 662 -258 663 -256
rect 665 -258 666 -256
rect 662 -259 666 -258
rect 929 -256 933 -241
rect 1112 -244 1116 -174
rect 1136 -95 1140 -94
rect 1371 -95 1375 -94
rect 1379 -29 1383 39
rect 1379 -31 1380 -29
rect 1382 -31 1383 -29
rect 1136 -97 1137 -95
rect 1139 -97 1140 -95
rect 1136 -184 1140 -97
rect 1379 -103 1383 -31
rect 1403 49 1407 50
rect 1638 49 1642 50
rect 1646 116 1650 183
rect 1646 114 1647 116
rect 1649 114 1650 116
rect 1403 47 1404 49
rect 1406 47 1407 49
rect 1403 -40 1407 47
rect 1646 41 1650 114
rect 1670 193 1674 194
rect 1670 191 1671 193
rect 1673 191 1674 193
rect 1670 104 1674 191
rect 1670 102 1671 104
rect 1673 102 1674 104
rect 1670 101 1674 102
rect 1686 129 1690 130
rect 1686 127 1687 129
rect 1689 127 1690 129
rect 1686 74 1690 127
rect 1686 72 1687 74
rect 1689 72 1690 74
rect 1686 71 1690 72
rect 1646 39 1647 41
rect 1649 39 1650 41
rect 1403 -42 1404 -40
rect 1406 -42 1407 -40
rect 1403 -43 1407 -42
rect 1419 -15 1423 -14
rect 1419 -17 1420 -15
rect 1422 -17 1423 -15
rect 1419 -70 1423 -17
rect 1419 -72 1420 -70
rect 1422 -72 1423 -70
rect 1419 -73 1423 -72
rect 1638 -27 1642 -26
rect 1638 -29 1639 -27
rect 1641 -29 1642 -27
rect 1638 -92 1642 -29
rect 1638 -94 1639 -92
rect 1641 -94 1642 -92
rect 1379 -105 1380 -103
rect 1382 -105 1383 -103
rect 1136 -186 1137 -184
rect 1139 -186 1140 -184
rect 1136 -187 1140 -186
rect 1152 -159 1156 -158
rect 1152 -161 1153 -159
rect 1155 -161 1156 -159
rect 1152 -214 1156 -161
rect 1152 -216 1153 -214
rect 1155 -216 1156 -214
rect 1152 -217 1156 -216
rect 1371 -171 1375 -170
rect 1371 -173 1372 -171
rect 1374 -173 1375 -171
rect 1371 -236 1375 -173
rect 1371 -238 1372 -236
rect 1374 -238 1375 -236
rect 1112 -246 1113 -244
rect 1115 -246 1116 -244
rect 1112 -247 1116 -246
rect 1196 -239 1200 -238
rect 1371 -239 1375 -238
rect 1379 -172 1383 -105
rect 1379 -174 1380 -172
rect 1382 -174 1383 -172
rect 1196 -241 1197 -239
rect 1199 -241 1200 -239
rect 929 -258 930 -256
rect 932 -258 933 -256
rect 929 -259 933 -258
rect 1196 -256 1200 -241
rect 1379 -244 1383 -174
rect 1403 -95 1407 -94
rect 1638 -95 1642 -94
rect 1646 -29 1650 39
rect 1646 -31 1647 -29
rect 1649 -31 1650 -29
rect 1403 -97 1404 -95
rect 1406 -97 1407 -95
rect 1403 -184 1407 -97
rect 1646 -103 1650 -31
rect 1670 49 1674 50
rect 1670 47 1671 49
rect 1673 47 1674 49
rect 1670 -40 1674 47
rect 1670 -42 1671 -40
rect 1673 -42 1674 -40
rect 1670 -43 1674 -42
rect 1686 -15 1690 -14
rect 1686 -17 1687 -15
rect 1689 -17 1690 -15
rect 1686 -70 1690 -17
rect 1686 -72 1687 -70
rect 1689 -72 1690 -70
rect 1686 -73 1690 -72
rect 1646 -105 1647 -103
rect 1649 -105 1650 -103
rect 1403 -186 1404 -184
rect 1406 -186 1407 -184
rect 1403 -187 1407 -186
rect 1419 -159 1423 -158
rect 1419 -161 1420 -159
rect 1422 -161 1423 -159
rect 1419 -214 1423 -161
rect 1419 -216 1420 -214
rect 1422 -216 1423 -214
rect 1419 -217 1423 -216
rect 1638 -171 1642 -170
rect 1638 -173 1639 -171
rect 1641 -173 1642 -171
rect 1638 -236 1642 -173
rect 1638 -238 1639 -236
rect 1641 -238 1642 -236
rect 1379 -246 1380 -244
rect 1382 -246 1383 -244
rect 1379 -247 1383 -246
rect 1463 -239 1467 -238
rect 1638 -239 1642 -238
rect 1646 -172 1650 -105
rect 1646 -174 1647 -172
rect 1649 -174 1650 -172
rect 1463 -241 1464 -239
rect 1466 -241 1467 -239
rect 1196 -258 1197 -256
rect 1199 -258 1200 -256
rect 1196 -259 1200 -258
rect 1463 -256 1467 -241
rect 1646 -244 1650 -174
rect 1670 -95 1674 -94
rect 1670 -97 1671 -95
rect 1673 -97 1674 -95
rect 1670 -184 1674 -97
rect 1670 -186 1671 -184
rect 1673 -186 1674 -184
rect 1670 -187 1674 -186
rect 1686 -159 1690 -158
rect 1686 -161 1687 -159
rect 1689 -161 1690 -159
rect 1686 -214 1690 -161
rect 1686 -216 1687 -214
rect 1689 -216 1690 -214
rect 1686 -217 1690 -216
rect 1769 -235 1773 300
rect 1928 290 1932 291
rect 1928 288 1929 290
rect 1931 288 1932 290
rect 1860 286 1864 287
rect 1860 284 1861 286
rect 1863 284 1864 286
rect 1814 273 1818 274
rect 1814 271 1815 273
rect 1817 271 1818 273
rect 1814 236 1818 271
rect 1860 273 1864 284
rect 1860 271 1861 273
rect 1863 271 1864 273
rect 1860 269 1864 271
rect 1814 234 1815 236
rect 1817 234 1818 236
rect 1814 233 1818 234
rect 1905 261 1909 262
rect 1905 259 1906 261
rect 1908 259 1909 261
rect 1880 218 1884 219
rect 1880 216 1881 218
rect 1883 216 1884 218
rect 1872 113 1876 114
rect 1872 111 1873 113
rect 1875 111 1876 113
rect 1864 79 1868 80
rect 1864 77 1865 79
rect 1867 77 1868 79
rect 1856 -32 1860 -31
rect 1856 -34 1857 -32
rect 1859 -34 1860 -32
rect 1848 -70 1852 -69
rect 1848 -72 1849 -70
rect 1851 -72 1852 -70
rect 1759 -236 1773 -235
rect 1759 -238 1760 -236
rect 1762 -238 1773 -236
rect 1646 -246 1647 -244
rect 1649 -246 1650 -244
rect 1646 -247 1650 -246
rect 1730 -239 1734 -238
rect 1759 -239 1773 -238
rect 1840 -176 1844 -175
rect 1840 -178 1841 -176
rect 1843 -178 1844 -176
rect 1730 -241 1731 -239
rect 1733 -241 1734 -239
rect 1463 -258 1464 -256
rect 1466 -258 1467 -256
rect 1463 -259 1467 -258
rect 1730 -256 1734 -241
rect 1840 -253 1844 -178
rect 1840 -255 1841 -253
rect 1843 -255 1844 -253
rect 1840 -256 1844 -255
rect 1730 -258 1731 -256
rect 1733 -258 1734 -256
rect 1730 -259 1734 -258
rect 1848 -261 1852 -72
rect 1848 -263 1849 -261
rect 1851 -263 1852 -261
rect 1848 -264 1852 -263
rect 1856 -269 1860 -34
rect 1864 -237 1868 77
rect 1864 -239 1865 -237
rect 1867 -239 1868 -237
rect 1864 -240 1868 -239
rect 1872 -245 1876 111
rect 1872 -247 1873 -245
rect 1875 -247 1876 -245
rect 1872 -248 1876 -247
rect 1880 -253 1884 216
rect 1905 196 1909 259
rect 1905 194 1906 196
rect 1908 194 1909 196
rect 1905 193 1909 194
rect 1928 256 1932 288
rect 2091 290 2095 291
rect 2091 288 2092 290
rect 2094 288 2095 290
rect 2091 273 2095 288
rect 2091 271 2092 273
rect 2094 271 2095 273
rect 2091 270 2095 271
rect 2192 273 2196 300
rect 2192 271 2193 273
rect 2195 271 2196 273
rect 2192 270 2196 271
rect 2263 303 2267 304
rect 2263 301 2264 303
rect 2266 301 2267 303
rect 1928 254 1929 256
rect 1931 254 1932 256
rect 1928 210 1932 254
rect 1928 208 1929 210
rect 1931 208 1932 210
rect 1905 117 1909 118
rect 1905 115 1906 117
rect 1908 115 1909 117
rect 1905 52 1909 115
rect 1905 50 1906 52
rect 1908 50 1909 52
rect 1905 49 1909 50
rect 1928 112 1932 208
rect 2191 261 2195 262
rect 2191 259 2192 261
rect 2194 259 2195 261
rect 2191 196 2195 259
rect 2263 235 2267 301
rect 2271 303 2275 304
rect 2271 301 2272 303
rect 2274 301 2275 303
rect 2271 243 2275 301
rect 2279 303 2283 304
rect 2279 301 2280 303
rect 2282 301 2283 303
rect 2279 251 2283 301
rect 2287 303 2291 304
rect 2287 301 2288 303
rect 2290 301 2291 303
rect 2287 259 2291 301
rect 2295 303 2299 304
rect 2295 301 2296 303
rect 2298 301 2299 303
rect 2295 267 2299 301
rect 2303 303 2307 304
rect 2303 301 2304 303
rect 2306 301 2307 303
rect 2303 274 2307 301
rect 2323 303 2331 304
rect 2323 301 2324 303
rect 2326 301 2328 303
rect 2330 301 2331 303
rect 2323 300 2331 301
rect 2303 272 2304 274
rect 2306 272 2307 274
rect 2303 271 2307 272
rect 2295 263 2307 267
rect 2287 255 2299 259
rect 2279 247 2291 251
rect 2271 239 2283 243
rect 2263 231 2275 235
rect 2263 226 2267 227
rect 2263 224 2264 226
rect 2266 224 2267 226
rect 2235 204 2239 205
rect 2235 202 2236 204
rect 2238 202 2239 204
rect 2235 200 2239 202
rect 2235 198 2236 200
rect 2238 198 2239 200
rect 2235 197 2239 198
rect 2191 194 2192 196
rect 2194 194 2195 196
rect 2191 193 2195 194
rect 2263 154 2267 224
rect 2271 162 2275 231
rect 2279 171 2283 239
rect 2287 179 2291 247
rect 2295 187 2299 255
rect 2303 194 2307 263
rect 2314 233 2318 234
rect 2314 231 2315 233
rect 2317 231 2318 233
rect 2314 229 2318 231
rect 2314 227 2315 229
rect 2317 227 2318 229
rect 2314 226 2318 227
rect 2303 192 2304 194
rect 2306 192 2307 194
rect 2303 191 2307 192
rect 2295 183 2307 187
rect 2287 175 2299 179
rect 2279 167 2291 171
rect 2271 158 2283 162
rect 2263 150 2275 154
rect 2227 137 2231 138
rect 2227 135 2228 137
rect 2230 135 2231 137
rect 2227 129 2231 135
rect 2227 127 2228 129
rect 2230 127 2231 129
rect 2227 126 2231 127
rect 1928 110 1929 112
rect 1931 110 1932 112
rect 1928 66 1932 110
rect 1928 64 1929 66
rect 1931 64 1932 66
rect 1905 -27 1909 -26
rect 1905 -29 1906 -27
rect 1908 -29 1909 -27
rect 1905 -92 1909 -29
rect 1905 -94 1906 -92
rect 1908 -94 1909 -92
rect 1905 -95 1909 -94
rect 1928 -32 1932 64
rect 2191 117 2195 118
rect 2191 115 2192 117
rect 2194 115 2195 117
rect 2191 52 2195 115
rect 2191 50 2192 52
rect 2194 50 2195 52
rect 2191 49 2195 50
rect 2219 67 2223 68
rect 2219 65 2220 67
rect 2222 65 2223 67
rect 2219 50 2223 65
rect 2219 48 2220 50
rect 2222 48 2223 50
rect 2219 47 2223 48
rect 2211 -17 2231 -16
rect 2211 -19 2212 -17
rect 2214 -19 2228 -17
rect 2230 -19 2231 -17
rect 2211 -20 2231 -19
rect 1928 -34 1929 -32
rect 1931 -34 1932 -32
rect 1928 -78 1932 -34
rect 1928 -80 1929 -78
rect 1931 -80 1932 -78
rect 1905 -171 1909 -170
rect 1905 -173 1906 -171
rect 1908 -173 1909 -171
rect 1880 -255 1881 -253
rect 1883 -255 1884 -253
rect 1880 -256 1884 -255
rect 1888 -214 1892 -213
rect 1888 -216 1889 -214
rect 1891 -216 1892 -214
rect 1888 -261 1892 -216
rect 1905 -236 1909 -173
rect 1928 -176 1932 -80
rect 2191 -27 2195 -26
rect 2191 -29 2192 -27
rect 2194 -29 2195 -27
rect 2191 -92 2195 -29
rect 2191 -94 2192 -92
rect 2194 -94 2195 -92
rect 2191 -95 2195 -94
rect 2203 -99 2239 -98
rect 2203 -101 2204 -99
rect 2206 -101 2236 -99
rect 2238 -101 2239 -99
rect 2203 -102 2239 -101
rect 2195 -154 2199 -153
rect 2195 -156 2196 -154
rect 2198 -156 2199 -154
rect 2195 -162 2199 -156
rect 2195 -164 2196 -162
rect 2198 -164 2199 -162
rect 2195 -165 2199 -164
rect 1928 -178 1929 -176
rect 1931 -178 1932 -176
rect 1928 -222 1932 -178
rect 1928 -224 1929 -222
rect 1931 -224 1932 -222
rect 1928 -225 1932 -224
rect 2191 -171 2195 -170
rect 2191 -173 2192 -171
rect 2194 -173 2195 -171
rect 1905 -238 1906 -236
rect 1908 -238 1909 -236
rect 1905 -239 1909 -238
rect 2191 -236 2195 -173
rect 2271 -198 2275 150
rect 2279 107 2283 158
rect 2287 115 2291 167
rect 2295 123 2299 175
rect 2303 130 2307 183
rect 2323 167 2331 168
rect 2323 165 2324 167
rect 2326 165 2328 167
rect 2330 165 2331 167
rect 2323 164 2331 165
rect 2303 128 2304 130
rect 2306 128 2307 130
rect 2303 127 2307 128
rect 2295 119 2307 123
rect 2287 111 2299 115
rect 2279 103 2291 107
rect 2287 35 2291 103
rect 2295 43 2299 111
rect 2303 50 2307 119
rect 2314 89 2318 90
rect 2314 87 2315 89
rect 2317 87 2318 89
rect 2314 85 2318 87
rect 2314 83 2315 85
rect 2317 83 2318 85
rect 2314 82 2318 83
rect 2303 48 2304 50
rect 2306 48 2307 50
rect 2303 47 2307 48
rect 2295 39 2307 43
rect 2287 31 2299 35
rect 2295 -21 2299 31
rect 2303 -14 2307 39
rect 2323 23 2331 24
rect 2323 21 2324 23
rect 2326 21 2328 23
rect 2330 21 2331 23
rect 2323 20 2331 21
rect 2303 -16 2304 -14
rect 2306 -16 2307 -14
rect 2303 -17 2307 -16
rect 2295 -25 2307 -21
rect 2303 -94 2307 -25
rect 2314 -55 2318 -54
rect 2314 -57 2315 -55
rect 2317 -57 2318 -55
rect 2314 -59 2318 -57
rect 2314 -61 2315 -59
rect 2317 -61 2318 -59
rect 2314 -62 2318 -61
rect 2303 -96 2304 -94
rect 2306 -96 2307 -94
rect 2303 -97 2307 -96
rect 2323 -121 2331 -120
rect 2323 -123 2324 -121
rect 2326 -123 2328 -121
rect 2330 -123 2331 -121
rect 2323 -124 2331 -123
rect 2307 -158 2315 -157
rect 2307 -160 2308 -158
rect 2310 -160 2312 -158
rect 2314 -160 2315 -158
rect 2307 -161 2315 -160
rect 2199 -202 2275 -198
rect 2327 -193 2331 -192
rect 2327 -195 2328 -193
rect 2330 -195 2331 -193
rect 2199 -228 2203 -202
rect 2327 -205 2331 -195
rect 2327 -207 2328 -205
rect 2330 -207 2331 -205
rect 2327 -208 2331 -207
rect 2199 -230 2200 -228
rect 2202 -230 2203 -228
rect 2199 -231 2203 -230
rect 2243 -227 2247 -226
rect 2243 -229 2244 -227
rect 2246 -229 2247 -227
rect 2191 -238 2192 -236
rect 2194 -238 2195 -236
rect 2191 -239 2195 -238
rect 2243 -240 2247 -229
rect 2243 -242 2244 -240
rect 2246 -242 2247 -240
rect 2243 -243 2247 -242
rect 2319 -238 2323 -237
rect 2319 -240 2320 -238
rect 2322 -240 2323 -238
rect 1888 -263 1889 -261
rect 1891 -263 1892 -261
rect 1888 -264 1892 -263
rect 1896 -256 1900 -255
rect 1896 -258 1897 -256
rect 1899 -258 1900 -256
rect 1856 -271 1857 -269
rect 1859 -271 1860 -269
rect 1856 -272 1860 -271
rect 1896 -268 1900 -258
rect 2319 -268 2323 -240
rect 1896 -272 2323 -268
rect 2327 -269 2337 -268
rect 2327 -271 2328 -269
rect 2330 -271 2334 -269
rect 2336 -271 2337 -269
rect 2327 -272 2337 -271
<< alu4 >>
rect 2263 303 2267 304
rect 2263 301 2264 303
rect 2266 301 2267 303
rect 2263 300 2267 301
rect 2271 303 2275 304
rect 2271 301 2272 303
rect 2274 301 2275 303
rect 2271 300 2275 301
rect 2279 303 2283 304
rect 2279 301 2280 303
rect 2282 301 2283 303
rect 2279 300 2283 301
rect 2287 303 2291 304
rect 2287 301 2288 303
rect 2290 301 2291 303
rect 1851 291 2239 295
rect 1851 287 1855 291
rect 262 286 1855 287
rect 262 284 263 286
rect 265 284 1855 286
rect 262 283 1855 284
rect 1860 286 1864 287
rect 1860 284 1861 286
rect 1863 284 1864 286
rect 1860 283 1864 284
rect 1869 283 2231 287
rect 1869 279 1873 283
rect 525 278 1873 279
rect 525 276 530 278
rect 532 276 1873 278
rect 525 275 1873 276
rect 1877 275 2223 279
rect 1877 271 1881 275
rect 796 270 1881 271
rect 796 268 797 270
rect 799 268 1881 270
rect 796 267 1881 268
rect 1885 267 2215 271
rect 1885 263 1889 267
rect 1063 262 1889 263
rect 1063 260 1064 262
rect 1066 260 1889 262
rect 1063 259 1889 260
rect 1893 259 2207 263
rect 1893 255 1897 259
rect 1330 254 1897 255
rect 1330 252 1331 254
rect 1333 252 1897 254
rect 1330 251 1897 252
rect 1901 251 2199 255
rect 1901 247 1905 251
rect 1597 246 1905 247
rect 1597 244 1598 246
rect 1600 244 1905 246
rect 1597 243 1905 244
rect 2195 -154 2199 251
rect 2203 -99 2207 259
rect 2211 -17 2215 267
rect 2219 67 2223 275
rect 2227 137 2231 283
rect 2235 204 2239 291
rect 2235 202 2236 204
rect 2238 202 2239 204
rect 2235 201 2239 202
rect 2243 282 2247 283
rect 2243 280 2244 282
rect 2246 280 2247 282
rect 2227 135 2228 137
rect 2230 135 2231 137
rect 2227 134 2231 135
rect 2219 65 2220 67
rect 2222 65 2223 67
rect 2219 64 2223 65
rect 2211 -19 2212 -17
rect 2214 -19 2215 -17
rect 2211 -20 2215 -19
rect 2203 -101 2204 -99
rect 2206 -101 2207 -99
rect 2203 -102 2207 -101
rect 2195 -156 2196 -154
rect 2198 -156 2199 -154
rect 2195 -157 2199 -156
rect 2243 -227 2247 280
rect 2243 -229 2244 -227
rect 2246 -229 2247 -227
rect 2243 -230 2247 -229
rect 36 -236 1763 -235
rect 2287 -236 2291 301
rect 36 -238 37 -236
rect 39 -238 1760 -236
rect 1762 -238 1763 -236
rect 36 -239 1763 -238
rect 1864 -237 2291 -236
rect 1864 -239 1865 -237
rect 1867 -239 2291 -237
rect 1864 -240 2291 -239
rect 2295 303 2299 304
rect 2295 301 2296 303
rect 2298 301 2299 303
rect 2295 -244 2299 301
rect 1872 -245 2299 -244
rect 1872 -247 1873 -245
rect 1875 -247 2299 -245
rect 1872 -248 2299 -247
rect 2303 303 2307 304
rect 2303 301 2304 303
rect 2306 301 2307 303
rect 2303 -252 2307 301
rect 2327 303 2337 304
rect 2327 301 2328 303
rect 2330 301 2334 303
rect 2336 301 2337 303
rect 2327 300 2337 301
rect 2314 233 2322 234
rect 2314 231 2315 233
rect 2317 231 2319 233
rect 2321 231 2322 233
rect 2314 230 2322 231
rect 2327 167 2337 168
rect 2327 165 2328 167
rect 2330 165 2334 167
rect 2336 165 2337 167
rect 2327 164 2337 165
rect 2314 89 2322 90
rect 2314 87 2315 89
rect 2317 87 2319 89
rect 2321 87 2322 89
rect 2314 86 2322 87
rect 2327 23 2337 24
rect 2327 21 2328 23
rect 2330 21 2334 23
rect 2336 21 2337 23
rect 2327 20 2337 21
rect 2314 -55 2322 -54
rect 2314 -57 2315 -55
rect 2317 -57 2319 -55
rect 2321 -57 2322 -55
rect 2314 -58 2322 -57
rect 2327 -121 2337 -120
rect 2327 -123 2328 -121
rect 2330 -123 2334 -121
rect 2336 -123 2337 -121
rect 2327 -124 2337 -123
rect 1840 -253 1852 -252
rect 1840 -255 1841 -253
rect 1843 -255 1849 -253
rect 1851 -255 1852 -253
rect 1840 -256 1852 -255
rect 1880 -253 2307 -252
rect 1880 -255 1881 -253
rect 1883 -255 2307 -253
rect 1880 -256 2307 -255
rect 2311 -158 2315 -157
rect 2311 -160 2312 -158
rect 2314 -160 2315 -158
rect 2311 -260 2315 -160
rect 2323 -205 2331 -204
rect 2323 -207 2324 -205
rect 2326 -207 2328 -205
rect 2330 -207 2331 -205
rect 2323 -208 2331 -207
rect 1848 -261 1860 -260
rect 1848 -263 1849 -261
rect 1851 -263 1857 -261
rect 1859 -263 1860 -261
rect 1848 -264 1860 -263
rect 1888 -261 2315 -260
rect 1888 -263 1889 -261
rect 1891 -263 2315 -261
rect 1888 -264 2315 -263
rect 2333 -265 2337 -264
rect 2333 -267 2334 -265
rect 2336 -267 2337 -265
rect 1856 -269 2283 -268
rect 1856 -271 1857 -269
rect 1859 -271 2280 -269
rect 2282 -271 2283 -269
rect 1856 -272 2283 -271
rect 2333 -269 2337 -267
rect 2333 -271 2334 -269
rect 2336 -271 2337 -269
rect 2333 -272 2337 -271
<< alu5 >>
rect -8 310 2341 318
rect -8 -278 0 310
rect 2263 303 2267 304
rect 2263 301 2264 303
rect 2266 301 2267 303
rect 1860 286 1864 287
rect 1860 284 1861 286
rect 1863 284 1864 286
rect 1860 283 1864 284
rect 1860 282 2247 283
rect 1860 280 2244 282
rect 2246 280 2247 282
rect 1860 279 2247 280
rect 2263 -252 2267 301
rect 1848 -253 2267 -252
rect 1848 -255 1849 -253
rect 1851 -255 2267 -253
rect 1848 -256 2267 -255
rect 2271 303 2275 304
rect 2271 301 2272 303
rect 2274 301 2275 303
rect 2271 -260 2275 301
rect 1856 -261 2275 -260
rect 1856 -263 1857 -261
rect 1859 -263 2275 -261
rect 1856 -264 2275 -263
rect 2279 303 2283 304
rect 2279 301 2280 303
rect 2282 301 2283 303
rect 2279 -269 2283 301
rect 2333 303 2341 310
rect 2333 301 2334 303
rect 2336 301 2341 303
rect 2319 234 2329 236
rect 2318 233 2323 234
rect 2318 231 2319 233
rect 2321 231 2323 233
rect 2318 230 2323 231
rect 2327 230 2329 234
rect 2319 228 2329 230
rect 2333 167 2341 301
rect 2333 165 2334 167
rect 2336 165 2341 167
rect 2319 90 2329 92
rect 2318 89 2323 90
rect 2318 87 2319 89
rect 2321 87 2323 89
rect 2318 86 2323 87
rect 2327 86 2329 90
rect 2319 84 2329 86
rect 2333 23 2341 165
rect 2333 21 2334 23
rect 2336 21 2341 23
rect 2319 -54 2329 -52
rect 2318 -55 2323 -54
rect 2318 -57 2319 -55
rect 2321 -57 2323 -55
rect 2318 -58 2323 -57
rect 2327 -58 2329 -54
rect 2319 -60 2329 -58
rect 2333 -121 2341 21
rect 2333 -123 2334 -121
rect 2336 -123 2341 -121
rect 2321 -198 2329 -196
rect 2321 -202 2323 -198
rect 2327 -202 2329 -198
rect 2321 -205 2329 -202
rect 2321 -207 2324 -205
rect 2326 -207 2329 -205
rect 2321 -208 2329 -207
rect 2279 -271 2280 -269
rect 2282 -271 2283 -269
rect 2279 -272 2283 -271
rect 2333 -265 2341 -123
rect 2333 -267 2334 -265
rect 2336 -267 2341 -265
rect 2333 -278 2341 -267
rect -8 -286 2341 -278
<< alu6 >>
rect -17 319 2350 327
rect -17 -287 -9 319
rect 2342 238 2350 319
rect 2319 234 2350 238
rect 2319 230 2323 234
rect 2327 230 2350 234
rect 2319 226 2350 230
rect 2342 94 2350 226
rect 2319 90 2350 94
rect 2319 86 2323 90
rect 2327 86 2350 90
rect 2319 82 2350 86
rect 2342 -50 2350 82
rect 2319 -54 2350 -50
rect 2319 -58 2323 -54
rect 2327 -58 2350 -54
rect 2319 -62 2350 -58
rect 2342 -194 2350 -62
rect 2319 -198 2350 -194
rect 2319 -202 2323 -198
rect 2327 -202 2350 -198
rect 2319 -206 2350 -202
rect 2342 -287 2350 -206
rect -17 -295 2350 -287
<< ptie >>
rect 37 239 43 241
rect 37 237 39 239
rect 41 237 43 239
rect 37 235 43 237
rect 77 239 83 241
rect 77 237 79 239
rect 81 237 83 239
rect 77 235 83 237
rect 296 239 302 241
rect 296 237 298 239
rect 300 237 302 239
rect 296 235 302 237
rect 344 239 350 241
rect 344 237 346 239
rect 348 237 350 239
rect 344 235 350 237
rect 563 239 569 241
rect 563 237 565 239
rect 567 237 569 239
rect 563 235 569 237
rect 611 239 617 241
rect 611 237 613 239
rect 615 237 617 239
rect 611 235 617 237
rect 830 239 836 241
rect 830 237 832 239
rect 834 237 836 239
rect 830 235 836 237
rect 878 239 884 241
rect 878 237 880 239
rect 882 237 884 239
rect 878 235 884 237
rect 1097 239 1103 241
rect 1097 237 1099 239
rect 1101 237 1103 239
rect 1097 235 1103 237
rect 1145 239 1151 241
rect 1145 237 1147 239
rect 1149 237 1151 239
rect 1145 235 1151 237
rect 1364 239 1370 241
rect 1364 237 1366 239
rect 1368 237 1370 239
rect 1364 235 1370 237
rect 1412 239 1418 241
rect 1412 237 1414 239
rect 1416 237 1418 239
rect 1412 235 1418 237
rect 1631 239 1637 241
rect 1631 237 1633 239
rect 1635 237 1637 239
rect 1631 235 1637 237
rect 1679 239 1685 241
rect 1679 237 1681 239
rect 1683 237 1685 239
rect 1679 235 1685 237
rect 1898 239 1904 241
rect 1898 237 1900 239
rect 1902 237 1904 239
rect 1898 235 1904 237
rect 1913 239 1919 241
rect 1913 237 1915 239
rect 1917 237 1919 239
rect 1913 235 1919 237
rect 2184 239 2190 241
rect 2184 237 2186 239
rect 2188 237 2190 239
rect 2184 235 2190 237
rect 37 227 43 229
rect 37 225 39 227
rect 41 225 43 227
rect 37 223 43 225
rect 77 227 83 229
rect 77 225 79 227
rect 81 225 83 227
rect 77 223 83 225
rect 296 227 302 229
rect 296 225 298 227
rect 300 225 302 227
rect 296 223 302 225
rect 344 227 350 229
rect 344 225 346 227
rect 348 225 350 227
rect 344 223 350 225
rect 563 227 569 229
rect 563 225 565 227
rect 567 225 569 227
rect 563 223 569 225
rect 611 227 617 229
rect 611 225 613 227
rect 615 225 617 227
rect 611 223 617 225
rect 830 227 836 229
rect 830 225 832 227
rect 834 225 836 227
rect 830 223 836 225
rect 878 227 884 229
rect 878 225 880 227
rect 882 225 884 227
rect 878 223 884 225
rect 1097 227 1103 229
rect 1097 225 1099 227
rect 1101 225 1103 227
rect 1097 223 1103 225
rect 1145 227 1151 229
rect 1145 225 1147 227
rect 1149 225 1151 227
rect 1145 223 1151 225
rect 1364 227 1370 229
rect 1364 225 1366 227
rect 1368 225 1370 227
rect 1364 223 1370 225
rect 1412 227 1418 229
rect 1412 225 1414 227
rect 1416 225 1418 227
rect 1412 223 1418 225
rect 1631 227 1637 229
rect 1631 225 1633 227
rect 1635 225 1637 227
rect 1631 223 1637 225
rect 1679 227 1685 229
rect 1679 225 1681 227
rect 1683 225 1685 227
rect 1679 223 1685 225
rect 1898 227 1904 229
rect 1898 225 1900 227
rect 1902 225 1904 227
rect 1898 223 1904 225
rect 1913 227 1919 229
rect 1913 225 1915 227
rect 1917 225 1919 227
rect 1913 223 1919 225
rect 2184 227 2190 229
rect 2184 225 2186 227
rect 2188 225 2190 227
rect 2184 223 2190 225
rect 37 95 43 97
rect 37 93 39 95
rect 41 93 43 95
rect 37 91 43 93
rect 77 95 83 97
rect 77 93 79 95
rect 81 93 83 95
rect 77 91 83 93
rect 296 95 302 97
rect 296 93 298 95
rect 300 93 302 95
rect 296 91 302 93
rect 344 95 350 97
rect 344 93 346 95
rect 348 93 350 95
rect 344 91 350 93
rect 563 95 569 97
rect 563 93 565 95
rect 567 93 569 95
rect 563 91 569 93
rect 611 95 617 97
rect 611 93 613 95
rect 615 93 617 95
rect 611 91 617 93
rect 830 95 836 97
rect 830 93 832 95
rect 834 93 836 95
rect 830 91 836 93
rect 878 95 884 97
rect 878 93 880 95
rect 882 93 884 95
rect 878 91 884 93
rect 1097 95 1103 97
rect 1097 93 1099 95
rect 1101 93 1103 95
rect 1097 91 1103 93
rect 1145 95 1151 97
rect 1145 93 1147 95
rect 1149 93 1151 95
rect 1145 91 1151 93
rect 1364 95 1370 97
rect 1364 93 1366 95
rect 1368 93 1370 95
rect 1364 91 1370 93
rect 1412 95 1418 97
rect 1412 93 1414 95
rect 1416 93 1418 95
rect 1412 91 1418 93
rect 1631 95 1637 97
rect 1631 93 1633 95
rect 1635 93 1637 95
rect 1631 91 1637 93
rect 1679 95 1685 97
rect 1679 93 1681 95
rect 1683 93 1685 95
rect 1679 91 1685 93
rect 1898 95 1904 97
rect 1898 93 1900 95
rect 1902 93 1904 95
rect 1898 91 1904 93
rect 1913 95 1919 97
rect 1913 93 1915 95
rect 1917 93 1919 95
rect 1913 91 1919 93
rect 2184 95 2190 97
rect 2184 93 2186 95
rect 2188 93 2190 95
rect 2184 91 2190 93
rect 37 83 43 85
rect 37 81 39 83
rect 41 81 43 83
rect 37 79 43 81
rect 77 83 83 85
rect 77 81 79 83
rect 81 81 83 83
rect 77 79 83 81
rect 296 83 302 85
rect 296 81 298 83
rect 300 81 302 83
rect 296 79 302 81
rect 344 83 350 85
rect 344 81 346 83
rect 348 81 350 83
rect 344 79 350 81
rect 563 83 569 85
rect 563 81 565 83
rect 567 81 569 83
rect 563 79 569 81
rect 611 83 617 85
rect 611 81 613 83
rect 615 81 617 83
rect 611 79 617 81
rect 830 83 836 85
rect 830 81 832 83
rect 834 81 836 83
rect 830 79 836 81
rect 878 83 884 85
rect 878 81 880 83
rect 882 81 884 83
rect 878 79 884 81
rect 1097 83 1103 85
rect 1097 81 1099 83
rect 1101 81 1103 83
rect 1097 79 1103 81
rect 1145 83 1151 85
rect 1145 81 1147 83
rect 1149 81 1151 83
rect 1145 79 1151 81
rect 1364 83 1370 85
rect 1364 81 1366 83
rect 1368 81 1370 83
rect 1364 79 1370 81
rect 1412 83 1418 85
rect 1412 81 1414 83
rect 1416 81 1418 83
rect 1412 79 1418 81
rect 1631 83 1637 85
rect 1631 81 1633 83
rect 1635 81 1637 83
rect 1631 79 1637 81
rect 1679 83 1685 85
rect 1679 81 1681 83
rect 1683 81 1685 83
rect 1679 79 1685 81
rect 1898 83 1904 85
rect 1898 81 1900 83
rect 1902 81 1904 83
rect 1898 79 1904 81
rect 1913 83 1919 85
rect 1913 81 1915 83
rect 1917 81 1919 83
rect 1913 79 1919 81
rect 2184 83 2190 85
rect 2184 81 2186 83
rect 2188 81 2190 83
rect 2184 79 2190 81
rect 37 -49 43 -47
rect 37 -51 39 -49
rect 41 -51 43 -49
rect 37 -53 43 -51
rect 77 -49 83 -47
rect 77 -51 79 -49
rect 81 -51 83 -49
rect 77 -53 83 -51
rect 296 -49 302 -47
rect 296 -51 298 -49
rect 300 -51 302 -49
rect 296 -53 302 -51
rect 344 -49 350 -47
rect 344 -51 346 -49
rect 348 -51 350 -49
rect 344 -53 350 -51
rect 563 -49 569 -47
rect 563 -51 565 -49
rect 567 -51 569 -49
rect 563 -53 569 -51
rect 611 -49 617 -47
rect 611 -51 613 -49
rect 615 -51 617 -49
rect 611 -53 617 -51
rect 830 -49 836 -47
rect 830 -51 832 -49
rect 834 -51 836 -49
rect 830 -53 836 -51
rect 878 -49 884 -47
rect 878 -51 880 -49
rect 882 -51 884 -49
rect 878 -53 884 -51
rect 1097 -49 1103 -47
rect 1097 -51 1099 -49
rect 1101 -51 1103 -49
rect 1097 -53 1103 -51
rect 1145 -49 1151 -47
rect 1145 -51 1147 -49
rect 1149 -51 1151 -49
rect 1145 -53 1151 -51
rect 1364 -49 1370 -47
rect 1364 -51 1366 -49
rect 1368 -51 1370 -49
rect 1364 -53 1370 -51
rect 1412 -49 1418 -47
rect 1412 -51 1414 -49
rect 1416 -51 1418 -49
rect 1412 -53 1418 -51
rect 1631 -49 1637 -47
rect 1631 -51 1633 -49
rect 1635 -51 1637 -49
rect 1631 -53 1637 -51
rect 1679 -49 1685 -47
rect 1679 -51 1681 -49
rect 1683 -51 1685 -49
rect 1679 -53 1685 -51
rect 1898 -49 1904 -47
rect 1898 -51 1900 -49
rect 1902 -51 1904 -49
rect 1898 -53 1904 -51
rect 1913 -49 1919 -47
rect 1913 -51 1915 -49
rect 1917 -51 1919 -49
rect 1913 -53 1919 -51
rect 2184 -49 2190 -47
rect 2184 -51 2186 -49
rect 2188 -51 2190 -49
rect 2184 -53 2190 -51
rect 37 -61 43 -59
rect 37 -63 39 -61
rect 41 -63 43 -61
rect 37 -65 43 -63
rect 77 -61 83 -59
rect 77 -63 79 -61
rect 81 -63 83 -61
rect 77 -65 83 -63
rect 296 -61 302 -59
rect 296 -63 298 -61
rect 300 -63 302 -61
rect 296 -65 302 -63
rect 344 -61 350 -59
rect 344 -63 346 -61
rect 348 -63 350 -61
rect 344 -65 350 -63
rect 563 -61 569 -59
rect 563 -63 565 -61
rect 567 -63 569 -61
rect 563 -65 569 -63
rect 611 -61 617 -59
rect 611 -63 613 -61
rect 615 -63 617 -61
rect 611 -65 617 -63
rect 830 -61 836 -59
rect 830 -63 832 -61
rect 834 -63 836 -61
rect 830 -65 836 -63
rect 878 -61 884 -59
rect 878 -63 880 -61
rect 882 -63 884 -61
rect 878 -65 884 -63
rect 1097 -61 1103 -59
rect 1097 -63 1099 -61
rect 1101 -63 1103 -61
rect 1097 -65 1103 -63
rect 1145 -61 1151 -59
rect 1145 -63 1147 -61
rect 1149 -63 1151 -61
rect 1145 -65 1151 -63
rect 1364 -61 1370 -59
rect 1364 -63 1366 -61
rect 1368 -63 1370 -61
rect 1364 -65 1370 -63
rect 1412 -61 1418 -59
rect 1412 -63 1414 -61
rect 1416 -63 1418 -61
rect 1412 -65 1418 -63
rect 1631 -61 1637 -59
rect 1631 -63 1633 -61
rect 1635 -63 1637 -61
rect 1631 -65 1637 -63
rect 1679 -61 1685 -59
rect 1679 -63 1681 -61
rect 1683 -63 1685 -61
rect 1679 -65 1685 -63
rect 1898 -61 1904 -59
rect 1898 -63 1900 -61
rect 1902 -63 1904 -61
rect 1898 -65 1904 -63
rect 1913 -61 1919 -59
rect 1913 -63 1915 -61
rect 1917 -63 1919 -61
rect 1913 -65 1919 -63
rect 2184 -61 2190 -59
rect 2184 -63 2186 -61
rect 2188 -63 2190 -61
rect 2184 -65 2190 -63
rect 37 -193 43 -191
rect 37 -195 39 -193
rect 41 -195 43 -193
rect 37 -197 43 -195
rect 77 -193 83 -191
rect 77 -195 79 -193
rect 81 -195 83 -193
rect 77 -197 83 -195
rect 296 -193 302 -191
rect 296 -195 298 -193
rect 300 -195 302 -193
rect 296 -197 302 -195
rect 344 -193 350 -191
rect 344 -195 346 -193
rect 348 -195 350 -193
rect 344 -197 350 -195
rect 563 -193 569 -191
rect 563 -195 565 -193
rect 567 -195 569 -193
rect 563 -197 569 -195
rect 611 -193 617 -191
rect 611 -195 613 -193
rect 615 -195 617 -193
rect 611 -197 617 -195
rect 830 -193 836 -191
rect 830 -195 832 -193
rect 834 -195 836 -193
rect 830 -197 836 -195
rect 878 -193 884 -191
rect 878 -195 880 -193
rect 882 -195 884 -193
rect 878 -197 884 -195
rect 1097 -193 1103 -191
rect 1097 -195 1099 -193
rect 1101 -195 1103 -193
rect 1097 -197 1103 -195
rect 1145 -193 1151 -191
rect 1145 -195 1147 -193
rect 1149 -195 1151 -193
rect 1145 -197 1151 -195
rect 1364 -193 1370 -191
rect 1364 -195 1366 -193
rect 1368 -195 1370 -193
rect 1364 -197 1370 -195
rect 1412 -193 1418 -191
rect 1412 -195 1414 -193
rect 1416 -195 1418 -193
rect 1412 -197 1418 -195
rect 1631 -193 1637 -191
rect 1631 -195 1633 -193
rect 1635 -195 1637 -193
rect 1631 -197 1637 -195
rect 1679 -193 1685 -191
rect 1679 -195 1681 -193
rect 1683 -195 1685 -193
rect 1679 -197 1685 -195
rect 1898 -193 1904 -191
rect 1898 -195 1900 -193
rect 1902 -195 1904 -193
rect 1898 -197 1904 -195
rect 1913 -193 1919 -191
rect 1913 -195 1915 -193
rect 1917 -195 1919 -193
rect 1913 -197 1919 -195
rect 2184 -193 2190 -191
rect 2184 -195 2186 -193
rect 2188 -195 2190 -193
rect 2184 -197 2190 -195
rect 37 -205 43 -203
rect 37 -207 39 -205
rect 41 -207 43 -205
rect 37 -209 43 -207
rect 77 -205 83 -203
rect 77 -207 79 -205
rect 81 -207 83 -205
rect 77 -209 83 -207
rect 296 -205 302 -203
rect 296 -207 298 -205
rect 300 -207 302 -205
rect 296 -209 302 -207
rect 344 -205 350 -203
rect 344 -207 346 -205
rect 348 -207 350 -205
rect 344 -209 350 -207
rect 563 -205 569 -203
rect 563 -207 565 -205
rect 567 -207 569 -205
rect 563 -209 569 -207
rect 611 -205 617 -203
rect 611 -207 613 -205
rect 615 -207 617 -205
rect 611 -209 617 -207
rect 830 -205 836 -203
rect 830 -207 832 -205
rect 834 -207 836 -205
rect 830 -209 836 -207
rect 878 -205 884 -203
rect 878 -207 880 -205
rect 882 -207 884 -205
rect 878 -209 884 -207
rect 1097 -205 1103 -203
rect 1097 -207 1099 -205
rect 1101 -207 1103 -205
rect 1097 -209 1103 -207
rect 1145 -205 1151 -203
rect 1145 -207 1147 -205
rect 1149 -207 1151 -205
rect 1145 -209 1151 -207
rect 1364 -205 1370 -203
rect 1364 -207 1366 -205
rect 1368 -207 1370 -205
rect 1364 -209 1370 -207
rect 1412 -205 1418 -203
rect 1412 -207 1414 -205
rect 1416 -207 1418 -205
rect 1412 -209 1418 -207
rect 1631 -205 1637 -203
rect 1631 -207 1633 -205
rect 1635 -207 1637 -205
rect 1631 -209 1637 -207
rect 1679 -205 1685 -203
rect 1679 -207 1681 -205
rect 1683 -207 1685 -205
rect 1679 -209 1685 -207
rect 1898 -205 1904 -203
rect 1898 -207 1900 -205
rect 1902 -207 1904 -205
rect 1898 -209 1904 -207
rect 1913 -205 1919 -203
rect 1913 -207 1915 -205
rect 1917 -207 1919 -205
rect 1913 -209 1919 -207
rect 2184 -205 2190 -203
rect 2184 -207 2186 -205
rect 2188 -207 2190 -205
rect 2184 -209 2190 -207
<< ntie >>
rect 37 299 43 301
rect 37 297 39 299
rect 41 297 43 299
rect 37 295 43 297
rect 77 299 83 301
rect 77 297 79 299
rect 81 297 83 299
rect 77 295 83 297
rect 296 299 302 301
rect 296 297 298 299
rect 300 297 302 299
rect 296 295 302 297
rect 344 299 350 301
rect 344 297 346 299
rect 348 297 350 299
rect 344 295 350 297
rect 563 299 569 301
rect 563 297 565 299
rect 567 297 569 299
rect 563 295 569 297
rect 611 299 617 301
rect 611 297 613 299
rect 615 297 617 299
rect 611 295 617 297
rect 830 299 836 301
rect 830 297 832 299
rect 834 297 836 299
rect 830 295 836 297
rect 878 299 884 301
rect 878 297 880 299
rect 882 297 884 299
rect 878 295 884 297
rect 1097 299 1103 301
rect 1097 297 1099 299
rect 1101 297 1103 299
rect 1097 295 1103 297
rect 1145 299 1151 301
rect 1145 297 1147 299
rect 1149 297 1151 299
rect 1145 295 1151 297
rect 1364 299 1370 301
rect 1364 297 1366 299
rect 1368 297 1370 299
rect 1364 295 1370 297
rect 1412 299 1418 301
rect 1412 297 1414 299
rect 1416 297 1418 299
rect 1412 295 1418 297
rect 1631 299 1637 301
rect 1631 297 1633 299
rect 1635 297 1637 299
rect 1631 295 1637 297
rect 1679 299 1685 301
rect 1679 297 1681 299
rect 1683 297 1685 299
rect 1679 295 1685 297
rect 1898 299 1904 301
rect 1898 297 1900 299
rect 1902 297 1904 299
rect 1946 299 1952 301
rect 1898 295 1904 297
rect 1946 297 1948 299
rect 1950 297 1952 299
rect 1946 295 1952 297
rect 2184 299 2190 301
rect 2184 297 2186 299
rect 2188 297 2190 299
rect 2184 295 2190 297
rect 37 167 43 169
rect 37 165 39 167
rect 41 165 43 167
rect 37 163 43 165
rect 77 167 83 169
rect 77 165 79 167
rect 81 165 83 167
rect 77 163 83 165
rect 296 167 302 169
rect 296 165 298 167
rect 300 165 302 167
rect 296 163 302 165
rect 344 167 350 169
rect 344 165 346 167
rect 348 165 350 167
rect 344 163 350 165
rect 563 167 569 169
rect 563 165 565 167
rect 567 165 569 167
rect 563 163 569 165
rect 611 167 617 169
rect 611 165 613 167
rect 615 165 617 167
rect 611 163 617 165
rect 830 167 836 169
rect 830 165 832 167
rect 834 165 836 167
rect 830 163 836 165
rect 878 167 884 169
rect 878 165 880 167
rect 882 165 884 167
rect 878 163 884 165
rect 1097 167 1103 169
rect 1097 165 1099 167
rect 1101 165 1103 167
rect 1097 163 1103 165
rect 1145 167 1151 169
rect 1145 165 1147 167
rect 1149 165 1151 167
rect 1145 163 1151 165
rect 1364 167 1370 169
rect 1364 165 1366 167
rect 1368 165 1370 167
rect 1364 163 1370 165
rect 1412 167 1418 169
rect 1412 165 1414 167
rect 1416 165 1418 167
rect 1412 163 1418 165
rect 1631 167 1637 169
rect 1631 165 1633 167
rect 1635 165 1637 167
rect 1631 163 1637 165
rect 1679 167 1685 169
rect 1679 165 1681 167
rect 1683 165 1685 167
rect 1679 163 1685 165
rect 1898 167 1904 169
rect 1898 165 1900 167
rect 1902 165 1904 167
rect 1946 167 1952 169
rect 1898 163 1904 165
rect 1946 165 1948 167
rect 1950 165 1952 167
rect 1946 163 1952 165
rect 2184 167 2190 169
rect 2184 165 2186 167
rect 2188 165 2190 167
rect 2184 163 2190 165
rect 37 155 43 157
rect 37 153 39 155
rect 41 153 43 155
rect 37 151 43 153
rect 77 155 83 157
rect 77 153 79 155
rect 81 153 83 155
rect 77 151 83 153
rect 296 155 302 157
rect 296 153 298 155
rect 300 153 302 155
rect 296 151 302 153
rect 344 155 350 157
rect 344 153 346 155
rect 348 153 350 155
rect 344 151 350 153
rect 563 155 569 157
rect 563 153 565 155
rect 567 153 569 155
rect 563 151 569 153
rect 611 155 617 157
rect 611 153 613 155
rect 615 153 617 155
rect 611 151 617 153
rect 830 155 836 157
rect 830 153 832 155
rect 834 153 836 155
rect 830 151 836 153
rect 878 155 884 157
rect 878 153 880 155
rect 882 153 884 155
rect 878 151 884 153
rect 1097 155 1103 157
rect 1097 153 1099 155
rect 1101 153 1103 155
rect 1097 151 1103 153
rect 1145 155 1151 157
rect 1145 153 1147 155
rect 1149 153 1151 155
rect 1145 151 1151 153
rect 1364 155 1370 157
rect 1364 153 1366 155
rect 1368 153 1370 155
rect 1364 151 1370 153
rect 1412 155 1418 157
rect 1412 153 1414 155
rect 1416 153 1418 155
rect 1412 151 1418 153
rect 1631 155 1637 157
rect 1631 153 1633 155
rect 1635 153 1637 155
rect 1631 151 1637 153
rect 1679 155 1685 157
rect 1679 153 1681 155
rect 1683 153 1685 155
rect 1679 151 1685 153
rect 1898 155 1904 157
rect 1898 153 1900 155
rect 1902 153 1904 155
rect 1946 155 1952 157
rect 1898 151 1904 153
rect 1946 153 1948 155
rect 1950 153 1952 155
rect 1946 151 1952 153
rect 2184 155 2190 157
rect 2184 153 2186 155
rect 2188 153 2190 155
rect 2184 151 2190 153
rect 37 23 43 25
rect 37 21 39 23
rect 41 21 43 23
rect 37 19 43 21
rect 77 23 83 25
rect 77 21 79 23
rect 81 21 83 23
rect 77 19 83 21
rect 296 23 302 25
rect 296 21 298 23
rect 300 21 302 23
rect 296 19 302 21
rect 344 23 350 25
rect 344 21 346 23
rect 348 21 350 23
rect 344 19 350 21
rect 563 23 569 25
rect 563 21 565 23
rect 567 21 569 23
rect 563 19 569 21
rect 611 23 617 25
rect 611 21 613 23
rect 615 21 617 23
rect 611 19 617 21
rect 830 23 836 25
rect 830 21 832 23
rect 834 21 836 23
rect 830 19 836 21
rect 878 23 884 25
rect 878 21 880 23
rect 882 21 884 23
rect 878 19 884 21
rect 1097 23 1103 25
rect 1097 21 1099 23
rect 1101 21 1103 23
rect 1097 19 1103 21
rect 1145 23 1151 25
rect 1145 21 1147 23
rect 1149 21 1151 23
rect 1145 19 1151 21
rect 1364 23 1370 25
rect 1364 21 1366 23
rect 1368 21 1370 23
rect 1364 19 1370 21
rect 1412 23 1418 25
rect 1412 21 1414 23
rect 1416 21 1418 23
rect 1412 19 1418 21
rect 1631 23 1637 25
rect 1631 21 1633 23
rect 1635 21 1637 23
rect 1631 19 1637 21
rect 1679 23 1685 25
rect 1679 21 1681 23
rect 1683 21 1685 23
rect 1679 19 1685 21
rect 1898 23 1904 25
rect 1898 21 1900 23
rect 1902 21 1904 23
rect 1946 23 1952 25
rect 1898 19 1904 21
rect 1946 21 1948 23
rect 1950 21 1952 23
rect 1946 19 1952 21
rect 2184 23 2190 25
rect 2184 21 2186 23
rect 2188 21 2190 23
rect 2184 19 2190 21
rect 37 11 43 13
rect 37 9 39 11
rect 41 9 43 11
rect 37 7 43 9
rect 77 11 83 13
rect 77 9 79 11
rect 81 9 83 11
rect 77 7 83 9
rect 296 11 302 13
rect 296 9 298 11
rect 300 9 302 11
rect 296 7 302 9
rect 344 11 350 13
rect 344 9 346 11
rect 348 9 350 11
rect 344 7 350 9
rect 563 11 569 13
rect 563 9 565 11
rect 567 9 569 11
rect 563 7 569 9
rect 611 11 617 13
rect 611 9 613 11
rect 615 9 617 11
rect 611 7 617 9
rect 830 11 836 13
rect 830 9 832 11
rect 834 9 836 11
rect 830 7 836 9
rect 878 11 884 13
rect 878 9 880 11
rect 882 9 884 11
rect 878 7 884 9
rect 1097 11 1103 13
rect 1097 9 1099 11
rect 1101 9 1103 11
rect 1097 7 1103 9
rect 1145 11 1151 13
rect 1145 9 1147 11
rect 1149 9 1151 11
rect 1145 7 1151 9
rect 1364 11 1370 13
rect 1364 9 1366 11
rect 1368 9 1370 11
rect 1364 7 1370 9
rect 1412 11 1418 13
rect 1412 9 1414 11
rect 1416 9 1418 11
rect 1412 7 1418 9
rect 1631 11 1637 13
rect 1631 9 1633 11
rect 1635 9 1637 11
rect 1631 7 1637 9
rect 1679 11 1685 13
rect 1679 9 1681 11
rect 1683 9 1685 11
rect 1679 7 1685 9
rect 1898 11 1904 13
rect 1898 9 1900 11
rect 1902 9 1904 11
rect 1946 11 1952 13
rect 1898 7 1904 9
rect 1946 9 1948 11
rect 1950 9 1952 11
rect 1946 7 1952 9
rect 2184 11 2190 13
rect 2184 9 2186 11
rect 2188 9 2190 11
rect 2184 7 2190 9
rect 37 -121 43 -119
rect 37 -123 39 -121
rect 41 -123 43 -121
rect 37 -125 43 -123
rect 77 -121 83 -119
rect 77 -123 79 -121
rect 81 -123 83 -121
rect 77 -125 83 -123
rect 296 -121 302 -119
rect 296 -123 298 -121
rect 300 -123 302 -121
rect 296 -125 302 -123
rect 344 -121 350 -119
rect 344 -123 346 -121
rect 348 -123 350 -121
rect 344 -125 350 -123
rect 563 -121 569 -119
rect 563 -123 565 -121
rect 567 -123 569 -121
rect 563 -125 569 -123
rect 611 -121 617 -119
rect 611 -123 613 -121
rect 615 -123 617 -121
rect 611 -125 617 -123
rect 830 -121 836 -119
rect 830 -123 832 -121
rect 834 -123 836 -121
rect 830 -125 836 -123
rect 878 -121 884 -119
rect 878 -123 880 -121
rect 882 -123 884 -121
rect 878 -125 884 -123
rect 1097 -121 1103 -119
rect 1097 -123 1099 -121
rect 1101 -123 1103 -121
rect 1097 -125 1103 -123
rect 1145 -121 1151 -119
rect 1145 -123 1147 -121
rect 1149 -123 1151 -121
rect 1145 -125 1151 -123
rect 1364 -121 1370 -119
rect 1364 -123 1366 -121
rect 1368 -123 1370 -121
rect 1364 -125 1370 -123
rect 1412 -121 1418 -119
rect 1412 -123 1414 -121
rect 1416 -123 1418 -121
rect 1412 -125 1418 -123
rect 1631 -121 1637 -119
rect 1631 -123 1633 -121
rect 1635 -123 1637 -121
rect 1631 -125 1637 -123
rect 1679 -121 1685 -119
rect 1679 -123 1681 -121
rect 1683 -123 1685 -121
rect 1679 -125 1685 -123
rect 1898 -121 1904 -119
rect 1898 -123 1900 -121
rect 1902 -123 1904 -121
rect 1946 -121 1952 -119
rect 1898 -125 1904 -123
rect 1946 -123 1948 -121
rect 1950 -123 1952 -121
rect 1946 -125 1952 -123
rect 2184 -121 2190 -119
rect 2184 -123 2186 -121
rect 2188 -123 2190 -121
rect 2184 -125 2190 -123
rect 37 -133 43 -131
rect 37 -135 39 -133
rect 41 -135 43 -133
rect 37 -137 43 -135
rect 77 -133 83 -131
rect 77 -135 79 -133
rect 81 -135 83 -133
rect 77 -137 83 -135
rect 296 -133 302 -131
rect 296 -135 298 -133
rect 300 -135 302 -133
rect 296 -137 302 -135
rect 344 -133 350 -131
rect 344 -135 346 -133
rect 348 -135 350 -133
rect 344 -137 350 -135
rect 563 -133 569 -131
rect 563 -135 565 -133
rect 567 -135 569 -133
rect 563 -137 569 -135
rect 611 -133 617 -131
rect 611 -135 613 -133
rect 615 -135 617 -133
rect 611 -137 617 -135
rect 830 -133 836 -131
rect 830 -135 832 -133
rect 834 -135 836 -133
rect 830 -137 836 -135
rect 878 -133 884 -131
rect 878 -135 880 -133
rect 882 -135 884 -133
rect 878 -137 884 -135
rect 1097 -133 1103 -131
rect 1097 -135 1099 -133
rect 1101 -135 1103 -133
rect 1097 -137 1103 -135
rect 1145 -133 1151 -131
rect 1145 -135 1147 -133
rect 1149 -135 1151 -133
rect 1145 -137 1151 -135
rect 1364 -133 1370 -131
rect 1364 -135 1366 -133
rect 1368 -135 1370 -133
rect 1364 -137 1370 -135
rect 1412 -133 1418 -131
rect 1412 -135 1414 -133
rect 1416 -135 1418 -133
rect 1412 -137 1418 -135
rect 1631 -133 1637 -131
rect 1631 -135 1633 -133
rect 1635 -135 1637 -133
rect 1631 -137 1637 -135
rect 1679 -133 1685 -131
rect 1679 -135 1681 -133
rect 1683 -135 1685 -133
rect 1679 -137 1685 -135
rect 1898 -133 1904 -131
rect 1898 -135 1900 -133
rect 1902 -135 1904 -133
rect 1946 -133 1952 -131
rect 1898 -137 1904 -135
rect 1946 -135 1948 -133
rect 1950 -135 1952 -133
rect 1946 -137 1952 -135
rect 2184 -133 2190 -131
rect 2184 -135 2186 -133
rect 2188 -135 2190 -133
rect 2184 -137 2190 -135
rect 37 -265 43 -263
rect 37 -267 39 -265
rect 41 -267 43 -265
rect 37 -269 43 -267
rect 77 -265 83 -263
rect 77 -267 79 -265
rect 81 -267 83 -265
rect 77 -269 83 -267
rect 296 -265 302 -263
rect 296 -267 298 -265
rect 300 -267 302 -265
rect 296 -269 302 -267
rect 344 -265 350 -263
rect 344 -267 346 -265
rect 348 -267 350 -265
rect 344 -269 350 -267
rect 563 -265 569 -263
rect 563 -267 565 -265
rect 567 -267 569 -265
rect 563 -269 569 -267
rect 611 -265 617 -263
rect 611 -267 613 -265
rect 615 -267 617 -265
rect 611 -269 617 -267
rect 830 -265 836 -263
rect 830 -267 832 -265
rect 834 -267 836 -265
rect 830 -269 836 -267
rect 878 -265 884 -263
rect 878 -267 880 -265
rect 882 -267 884 -265
rect 878 -269 884 -267
rect 1097 -265 1103 -263
rect 1097 -267 1099 -265
rect 1101 -267 1103 -265
rect 1097 -269 1103 -267
rect 1145 -265 1151 -263
rect 1145 -267 1147 -265
rect 1149 -267 1151 -265
rect 1145 -269 1151 -267
rect 1364 -265 1370 -263
rect 1364 -267 1366 -265
rect 1368 -267 1370 -265
rect 1364 -269 1370 -267
rect 1412 -265 1418 -263
rect 1412 -267 1414 -265
rect 1416 -267 1418 -265
rect 1412 -269 1418 -267
rect 1631 -265 1637 -263
rect 1631 -267 1633 -265
rect 1635 -267 1637 -265
rect 1631 -269 1637 -267
rect 1679 -265 1685 -263
rect 1679 -267 1681 -265
rect 1683 -267 1685 -265
rect 1679 -269 1685 -267
rect 1898 -265 1904 -263
rect 1898 -267 1900 -265
rect 1902 -267 1904 -265
rect 1946 -265 1952 -263
rect 1898 -269 1904 -267
rect 1946 -267 1948 -265
rect 1950 -267 1952 -265
rect 1946 -269 1952 -267
rect 2184 -265 2190 -263
rect 2184 -267 2186 -265
rect 2188 -267 2190 -265
rect 2184 -269 2190 -267
<< nmos >>
rect 15 245 17 256
rect 22 245 24 256
rect 35 247 37 256
rect 55 245 57 256
rect 62 245 64 256
rect 75 247 77 256
rect 95 238 97 251
rect 105 241 107 251
rect 115 244 117 258
rect 125 244 127 258
rect 145 238 147 258
rect 152 238 154 258
rect 163 238 165 252
rect 185 238 187 252
rect 196 238 198 258
rect 203 238 205 258
rect 223 244 225 258
rect 233 244 235 258
rect 274 252 276 258
rect 284 252 286 258
rect 243 241 245 251
rect 253 238 255 251
rect 294 249 296 258
rect 322 245 324 256
rect 329 245 331 256
rect 342 247 344 256
rect 362 238 364 251
rect 372 241 374 251
rect 382 244 384 258
rect 392 244 394 258
rect 412 238 414 258
rect 419 238 421 258
rect 430 238 432 252
rect 452 238 454 252
rect 463 238 465 258
rect 470 238 472 258
rect 490 244 492 258
rect 500 244 502 258
rect 541 252 543 258
rect 551 252 553 258
rect 510 241 512 251
rect 520 238 522 251
rect 561 249 563 258
rect 589 245 591 256
rect 596 245 598 256
rect 609 247 611 256
rect 629 238 631 251
rect 639 241 641 251
rect 649 244 651 258
rect 659 244 661 258
rect 679 238 681 258
rect 686 238 688 258
rect 697 238 699 252
rect 719 238 721 252
rect 730 238 732 258
rect 737 238 739 258
rect 757 244 759 258
rect 767 244 769 258
rect 808 252 810 258
rect 818 252 820 258
rect 777 241 779 251
rect 787 238 789 251
rect 828 249 830 258
rect 856 245 858 256
rect 863 245 865 256
rect 876 247 878 256
rect 896 238 898 251
rect 906 241 908 251
rect 916 244 918 258
rect 926 244 928 258
rect 946 238 948 258
rect 953 238 955 258
rect 964 238 966 252
rect 986 238 988 252
rect 997 238 999 258
rect 1004 238 1006 258
rect 1024 244 1026 258
rect 1034 244 1036 258
rect 1075 252 1077 258
rect 1085 252 1087 258
rect 1044 241 1046 251
rect 1054 238 1056 251
rect 1095 249 1097 258
rect 1123 245 1125 256
rect 1130 245 1132 256
rect 1143 247 1145 256
rect 1163 238 1165 251
rect 1173 241 1175 251
rect 1183 244 1185 258
rect 1193 244 1195 258
rect 1213 238 1215 258
rect 1220 238 1222 258
rect 1231 238 1233 252
rect 1253 238 1255 252
rect 1264 238 1266 258
rect 1271 238 1273 258
rect 1291 244 1293 258
rect 1301 244 1303 258
rect 1342 252 1344 258
rect 1352 252 1354 258
rect 1311 241 1313 251
rect 1321 238 1323 251
rect 1362 249 1364 258
rect 1390 245 1392 256
rect 1397 245 1399 256
rect 1410 247 1412 256
rect 1430 238 1432 251
rect 1440 241 1442 251
rect 1450 244 1452 258
rect 1460 244 1462 258
rect 1480 238 1482 258
rect 1487 238 1489 258
rect 1498 238 1500 252
rect 1520 238 1522 252
rect 1531 238 1533 258
rect 1538 238 1540 258
rect 1558 244 1560 258
rect 1568 244 1570 258
rect 1609 252 1611 258
rect 1619 252 1621 258
rect 1578 241 1580 251
rect 1588 238 1590 251
rect 1629 249 1631 258
rect 1657 245 1659 256
rect 1664 245 1666 256
rect 1677 247 1679 256
rect 1697 238 1699 251
rect 1707 241 1709 251
rect 1717 244 1719 258
rect 1727 244 1729 258
rect 1747 238 1749 258
rect 1754 238 1756 258
rect 1765 238 1767 252
rect 1787 238 1789 252
rect 1798 238 1800 258
rect 1805 238 1807 258
rect 1825 244 1827 258
rect 1835 244 1837 258
rect 1876 252 1878 258
rect 1886 252 1888 258
rect 1845 241 1847 251
rect 1855 238 1857 251
rect 1896 249 1898 258
rect 1919 249 1921 258
rect 1935 244 1937 253
rect 1945 244 1947 253
rect 1955 241 1957 253
rect 1962 241 1964 253
rect 1983 238 1985 251
rect 1993 241 1995 251
rect 2003 244 2005 258
rect 2013 244 2015 258
rect 2033 238 2035 258
rect 2040 238 2042 258
rect 2051 238 2053 252
rect 2073 238 2075 252
rect 2084 238 2086 258
rect 2091 238 2093 258
rect 2111 244 2113 258
rect 2121 244 2123 258
rect 2162 252 2164 258
rect 2172 252 2174 258
rect 2131 241 2133 251
rect 2141 238 2143 251
rect 2182 249 2184 258
rect 2206 246 2208 252
rect 2216 244 2218 252
rect 2223 244 2225 252
rect 2233 244 2235 252
rect 2240 244 2242 252
rect 2250 244 2252 253
rect 2274 246 2276 252
rect 2284 244 2286 252
rect 2291 244 2293 252
rect 2301 244 2303 252
rect 2308 244 2310 252
rect 2318 244 2320 253
rect 15 208 17 219
rect 22 208 24 219
rect 35 208 37 217
rect 55 208 57 219
rect 62 208 64 219
rect 75 208 77 217
rect 95 213 97 226
rect 105 213 107 223
rect 115 206 117 220
rect 125 206 127 220
rect 145 206 147 226
rect 152 206 154 226
rect 163 212 165 226
rect 185 212 187 226
rect 196 206 198 226
rect 203 206 205 226
rect 223 206 225 220
rect 233 206 235 220
rect 243 213 245 223
rect 253 213 255 226
rect 274 206 276 212
rect 284 206 286 212
rect 294 206 296 215
rect 322 208 324 219
rect 329 208 331 219
rect 342 208 344 217
rect 362 213 364 226
rect 372 213 374 223
rect 382 206 384 220
rect 392 206 394 220
rect 412 206 414 226
rect 419 206 421 226
rect 430 212 432 226
rect 452 212 454 226
rect 463 206 465 226
rect 470 206 472 226
rect 490 206 492 220
rect 500 206 502 220
rect 510 213 512 223
rect 520 213 522 226
rect 541 206 543 212
rect 551 206 553 212
rect 561 206 563 215
rect 589 208 591 219
rect 596 208 598 219
rect 609 208 611 217
rect 629 213 631 226
rect 639 213 641 223
rect 649 206 651 220
rect 659 206 661 220
rect 679 206 681 226
rect 686 206 688 226
rect 697 212 699 226
rect 719 212 721 226
rect 730 206 732 226
rect 737 206 739 226
rect 757 206 759 220
rect 767 206 769 220
rect 777 213 779 223
rect 787 213 789 226
rect 808 206 810 212
rect 818 206 820 212
rect 828 206 830 215
rect 856 208 858 219
rect 863 208 865 219
rect 876 208 878 217
rect 896 213 898 226
rect 906 213 908 223
rect 916 206 918 220
rect 926 206 928 220
rect 946 206 948 226
rect 953 206 955 226
rect 964 212 966 226
rect 986 212 988 226
rect 997 206 999 226
rect 1004 206 1006 226
rect 1024 206 1026 220
rect 1034 206 1036 220
rect 1044 213 1046 223
rect 1054 213 1056 226
rect 1075 206 1077 212
rect 1085 206 1087 212
rect 1095 206 1097 215
rect 1123 208 1125 219
rect 1130 208 1132 219
rect 1143 208 1145 217
rect 1163 213 1165 226
rect 1173 213 1175 223
rect 1183 206 1185 220
rect 1193 206 1195 220
rect 1213 206 1215 226
rect 1220 206 1222 226
rect 1231 212 1233 226
rect 1253 212 1255 226
rect 1264 206 1266 226
rect 1271 206 1273 226
rect 1291 206 1293 220
rect 1301 206 1303 220
rect 1311 213 1313 223
rect 1321 213 1323 226
rect 1342 206 1344 212
rect 1352 206 1354 212
rect 1362 206 1364 215
rect 1390 208 1392 219
rect 1397 208 1399 219
rect 1410 208 1412 217
rect 1430 213 1432 226
rect 1440 213 1442 223
rect 1450 206 1452 220
rect 1460 206 1462 220
rect 1480 206 1482 226
rect 1487 206 1489 226
rect 1498 212 1500 226
rect 1520 212 1522 226
rect 1531 206 1533 226
rect 1538 206 1540 226
rect 1558 206 1560 220
rect 1568 206 1570 220
rect 1578 213 1580 223
rect 1588 213 1590 226
rect 1609 206 1611 212
rect 1619 206 1621 212
rect 1629 206 1631 215
rect 1657 208 1659 219
rect 1664 208 1666 219
rect 1677 208 1679 217
rect 1697 213 1699 226
rect 1707 213 1709 223
rect 1717 206 1719 220
rect 1727 206 1729 220
rect 1747 206 1749 226
rect 1754 206 1756 226
rect 1765 212 1767 226
rect 1787 212 1789 226
rect 1798 206 1800 226
rect 1805 206 1807 226
rect 1825 206 1827 220
rect 1835 206 1837 220
rect 1845 213 1847 223
rect 1855 213 1857 226
rect 1876 206 1878 212
rect 1886 206 1888 212
rect 1896 206 1898 215
rect 1919 206 1921 215
rect 1935 211 1937 220
rect 1945 211 1947 220
rect 1955 211 1957 223
rect 1962 211 1964 223
rect 1983 213 1985 226
rect 1993 213 1995 223
rect 2003 206 2005 220
rect 2013 206 2015 220
rect 2033 206 2035 226
rect 2040 206 2042 226
rect 2051 212 2053 226
rect 2073 212 2075 226
rect 2084 206 2086 226
rect 2091 206 2093 226
rect 2111 206 2113 220
rect 2121 206 2123 220
rect 2131 213 2133 223
rect 2141 213 2143 226
rect 2162 206 2164 212
rect 2172 206 2174 212
rect 2182 206 2184 215
rect 2206 212 2208 218
rect 2216 212 2218 220
rect 2223 212 2225 220
rect 2233 212 2235 220
rect 2240 212 2242 220
rect 2250 211 2252 220
rect 2274 212 2276 218
rect 2284 212 2286 220
rect 2291 212 2293 220
rect 2301 212 2303 220
rect 2308 212 2310 220
rect 2318 211 2320 220
rect 15 101 17 112
rect 22 101 24 112
rect 35 103 37 112
rect 55 101 57 112
rect 62 101 64 112
rect 75 103 77 112
rect 95 94 97 107
rect 105 97 107 107
rect 115 100 117 114
rect 125 100 127 114
rect 145 94 147 114
rect 152 94 154 114
rect 163 94 165 108
rect 185 94 187 108
rect 196 94 198 114
rect 203 94 205 114
rect 223 100 225 114
rect 233 100 235 114
rect 274 108 276 114
rect 284 108 286 114
rect 243 97 245 107
rect 253 94 255 107
rect 294 105 296 114
rect 322 101 324 112
rect 329 101 331 112
rect 342 103 344 112
rect 362 94 364 107
rect 372 97 374 107
rect 382 100 384 114
rect 392 100 394 114
rect 412 94 414 114
rect 419 94 421 114
rect 430 94 432 108
rect 452 94 454 108
rect 463 94 465 114
rect 470 94 472 114
rect 490 100 492 114
rect 500 100 502 114
rect 541 108 543 114
rect 551 108 553 114
rect 510 97 512 107
rect 520 94 522 107
rect 561 105 563 114
rect 589 101 591 112
rect 596 101 598 112
rect 609 103 611 112
rect 629 94 631 107
rect 639 97 641 107
rect 649 100 651 114
rect 659 100 661 114
rect 679 94 681 114
rect 686 94 688 114
rect 697 94 699 108
rect 719 94 721 108
rect 730 94 732 114
rect 737 94 739 114
rect 757 100 759 114
rect 767 100 769 114
rect 808 108 810 114
rect 818 108 820 114
rect 777 97 779 107
rect 787 94 789 107
rect 828 105 830 114
rect 856 101 858 112
rect 863 101 865 112
rect 876 103 878 112
rect 896 94 898 107
rect 906 97 908 107
rect 916 100 918 114
rect 926 100 928 114
rect 946 94 948 114
rect 953 94 955 114
rect 964 94 966 108
rect 986 94 988 108
rect 997 94 999 114
rect 1004 94 1006 114
rect 1024 100 1026 114
rect 1034 100 1036 114
rect 1075 108 1077 114
rect 1085 108 1087 114
rect 1044 97 1046 107
rect 1054 94 1056 107
rect 1095 105 1097 114
rect 1123 101 1125 112
rect 1130 101 1132 112
rect 1143 103 1145 112
rect 1163 94 1165 107
rect 1173 97 1175 107
rect 1183 100 1185 114
rect 1193 100 1195 114
rect 1213 94 1215 114
rect 1220 94 1222 114
rect 1231 94 1233 108
rect 1253 94 1255 108
rect 1264 94 1266 114
rect 1271 94 1273 114
rect 1291 100 1293 114
rect 1301 100 1303 114
rect 1342 108 1344 114
rect 1352 108 1354 114
rect 1311 97 1313 107
rect 1321 94 1323 107
rect 1362 105 1364 114
rect 1390 101 1392 112
rect 1397 101 1399 112
rect 1410 103 1412 112
rect 1430 94 1432 107
rect 1440 97 1442 107
rect 1450 100 1452 114
rect 1460 100 1462 114
rect 1480 94 1482 114
rect 1487 94 1489 114
rect 1498 94 1500 108
rect 1520 94 1522 108
rect 1531 94 1533 114
rect 1538 94 1540 114
rect 1558 100 1560 114
rect 1568 100 1570 114
rect 1609 108 1611 114
rect 1619 108 1621 114
rect 1578 97 1580 107
rect 1588 94 1590 107
rect 1629 105 1631 114
rect 1657 101 1659 112
rect 1664 101 1666 112
rect 1677 103 1679 112
rect 1697 94 1699 107
rect 1707 97 1709 107
rect 1717 100 1719 114
rect 1727 100 1729 114
rect 1747 94 1749 114
rect 1754 94 1756 114
rect 1765 94 1767 108
rect 1787 94 1789 108
rect 1798 94 1800 114
rect 1805 94 1807 114
rect 1825 100 1827 114
rect 1835 100 1837 114
rect 1876 108 1878 114
rect 1886 108 1888 114
rect 1845 97 1847 107
rect 1855 94 1857 107
rect 1896 105 1898 114
rect 1919 105 1921 114
rect 1935 100 1937 109
rect 1945 100 1947 109
rect 1955 97 1957 109
rect 1962 97 1964 109
rect 1983 94 1985 107
rect 1993 97 1995 107
rect 2003 100 2005 114
rect 2013 100 2015 114
rect 2033 94 2035 114
rect 2040 94 2042 114
rect 2051 94 2053 108
rect 2073 94 2075 108
rect 2084 94 2086 114
rect 2091 94 2093 114
rect 2111 100 2113 114
rect 2121 100 2123 114
rect 2162 108 2164 114
rect 2172 108 2174 114
rect 2131 97 2133 107
rect 2141 94 2143 107
rect 2182 105 2184 114
rect 2206 102 2208 108
rect 2216 100 2218 108
rect 2223 100 2225 108
rect 2233 100 2235 108
rect 2240 100 2242 108
rect 2250 100 2252 109
rect 2274 102 2276 108
rect 2284 100 2286 108
rect 2291 100 2293 108
rect 2301 100 2303 108
rect 2308 100 2310 108
rect 2318 100 2320 109
rect 15 64 17 75
rect 22 64 24 75
rect 35 64 37 73
rect 55 64 57 75
rect 62 64 64 75
rect 75 64 77 73
rect 95 69 97 82
rect 105 69 107 79
rect 115 62 117 76
rect 125 62 127 76
rect 145 62 147 82
rect 152 62 154 82
rect 163 68 165 82
rect 185 68 187 82
rect 196 62 198 82
rect 203 62 205 82
rect 223 62 225 76
rect 233 62 235 76
rect 243 69 245 79
rect 253 69 255 82
rect 274 62 276 68
rect 284 62 286 68
rect 294 62 296 71
rect 322 64 324 75
rect 329 64 331 75
rect 342 64 344 73
rect 362 69 364 82
rect 372 69 374 79
rect 382 62 384 76
rect 392 62 394 76
rect 412 62 414 82
rect 419 62 421 82
rect 430 68 432 82
rect 452 68 454 82
rect 463 62 465 82
rect 470 62 472 82
rect 490 62 492 76
rect 500 62 502 76
rect 510 69 512 79
rect 520 69 522 82
rect 541 62 543 68
rect 551 62 553 68
rect 561 62 563 71
rect 589 64 591 75
rect 596 64 598 75
rect 609 64 611 73
rect 629 69 631 82
rect 639 69 641 79
rect 649 62 651 76
rect 659 62 661 76
rect 679 62 681 82
rect 686 62 688 82
rect 697 68 699 82
rect 719 68 721 82
rect 730 62 732 82
rect 737 62 739 82
rect 757 62 759 76
rect 767 62 769 76
rect 777 69 779 79
rect 787 69 789 82
rect 808 62 810 68
rect 818 62 820 68
rect 828 62 830 71
rect 856 64 858 75
rect 863 64 865 75
rect 876 64 878 73
rect 896 69 898 82
rect 906 69 908 79
rect 916 62 918 76
rect 926 62 928 76
rect 946 62 948 82
rect 953 62 955 82
rect 964 68 966 82
rect 986 68 988 82
rect 997 62 999 82
rect 1004 62 1006 82
rect 1024 62 1026 76
rect 1034 62 1036 76
rect 1044 69 1046 79
rect 1054 69 1056 82
rect 1075 62 1077 68
rect 1085 62 1087 68
rect 1095 62 1097 71
rect 1123 64 1125 75
rect 1130 64 1132 75
rect 1143 64 1145 73
rect 1163 69 1165 82
rect 1173 69 1175 79
rect 1183 62 1185 76
rect 1193 62 1195 76
rect 1213 62 1215 82
rect 1220 62 1222 82
rect 1231 68 1233 82
rect 1253 68 1255 82
rect 1264 62 1266 82
rect 1271 62 1273 82
rect 1291 62 1293 76
rect 1301 62 1303 76
rect 1311 69 1313 79
rect 1321 69 1323 82
rect 1342 62 1344 68
rect 1352 62 1354 68
rect 1362 62 1364 71
rect 1390 64 1392 75
rect 1397 64 1399 75
rect 1410 64 1412 73
rect 1430 69 1432 82
rect 1440 69 1442 79
rect 1450 62 1452 76
rect 1460 62 1462 76
rect 1480 62 1482 82
rect 1487 62 1489 82
rect 1498 68 1500 82
rect 1520 68 1522 82
rect 1531 62 1533 82
rect 1538 62 1540 82
rect 1558 62 1560 76
rect 1568 62 1570 76
rect 1578 69 1580 79
rect 1588 69 1590 82
rect 1609 62 1611 68
rect 1619 62 1621 68
rect 1629 62 1631 71
rect 1657 64 1659 75
rect 1664 64 1666 75
rect 1677 64 1679 73
rect 1697 69 1699 82
rect 1707 69 1709 79
rect 1717 62 1719 76
rect 1727 62 1729 76
rect 1747 62 1749 82
rect 1754 62 1756 82
rect 1765 68 1767 82
rect 1787 68 1789 82
rect 1798 62 1800 82
rect 1805 62 1807 82
rect 1825 62 1827 76
rect 1835 62 1837 76
rect 1845 69 1847 79
rect 1855 69 1857 82
rect 1876 62 1878 68
rect 1886 62 1888 68
rect 1896 62 1898 71
rect 1919 62 1921 71
rect 1935 67 1937 76
rect 1945 67 1947 76
rect 1955 67 1957 79
rect 1962 67 1964 79
rect 1983 69 1985 82
rect 1993 69 1995 79
rect 2003 62 2005 76
rect 2013 62 2015 76
rect 2033 62 2035 82
rect 2040 62 2042 82
rect 2051 68 2053 82
rect 2073 68 2075 82
rect 2084 62 2086 82
rect 2091 62 2093 82
rect 2111 62 2113 76
rect 2121 62 2123 76
rect 2131 69 2133 79
rect 2141 69 2143 82
rect 2162 62 2164 68
rect 2172 62 2174 68
rect 2182 62 2184 71
rect 2206 68 2208 74
rect 2216 68 2218 76
rect 2223 68 2225 76
rect 2233 68 2235 76
rect 2240 68 2242 76
rect 2250 67 2252 76
rect 2274 68 2276 74
rect 2284 68 2286 76
rect 2291 68 2293 76
rect 2301 68 2303 76
rect 2308 68 2310 76
rect 2318 67 2320 76
rect 15 -43 17 -32
rect 22 -43 24 -32
rect 35 -41 37 -32
rect 55 -43 57 -32
rect 62 -43 64 -32
rect 75 -41 77 -32
rect 95 -50 97 -37
rect 105 -47 107 -37
rect 115 -44 117 -30
rect 125 -44 127 -30
rect 145 -50 147 -30
rect 152 -50 154 -30
rect 163 -50 165 -36
rect 185 -50 187 -36
rect 196 -50 198 -30
rect 203 -50 205 -30
rect 223 -44 225 -30
rect 233 -44 235 -30
rect 274 -36 276 -30
rect 284 -36 286 -30
rect 243 -47 245 -37
rect 253 -50 255 -37
rect 294 -39 296 -30
rect 322 -43 324 -32
rect 329 -43 331 -32
rect 342 -41 344 -32
rect 362 -50 364 -37
rect 372 -47 374 -37
rect 382 -44 384 -30
rect 392 -44 394 -30
rect 412 -50 414 -30
rect 419 -50 421 -30
rect 430 -50 432 -36
rect 452 -50 454 -36
rect 463 -50 465 -30
rect 470 -50 472 -30
rect 490 -44 492 -30
rect 500 -44 502 -30
rect 541 -36 543 -30
rect 551 -36 553 -30
rect 510 -47 512 -37
rect 520 -50 522 -37
rect 561 -39 563 -30
rect 589 -43 591 -32
rect 596 -43 598 -32
rect 609 -41 611 -32
rect 629 -50 631 -37
rect 639 -47 641 -37
rect 649 -44 651 -30
rect 659 -44 661 -30
rect 679 -50 681 -30
rect 686 -50 688 -30
rect 697 -50 699 -36
rect 719 -50 721 -36
rect 730 -50 732 -30
rect 737 -50 739 -30
rect 757 -44 759 -30
rect 767 -44 769 -30
rect 808 -36 810 -30
rect 818 -36 820 -30
rect 777 -47 779 -37
rect 787 -50 789 -37
rect 828 -39 830 -30
rect 856 -43 858 -32
rect 863 -43 865 -32
rect 876 -41 878 -32
rect 896 -50 898 -37
rect 906 -47 908 -37
rect 916 -44 918 -30
rect 926 -44 928 -30
rect 946 -50 948 -30
rect 953 -50 955 -30
rect 964 -50 966 -36
rect 986 -50 988 -36
rect 997 -50 999 -30
rect 1004 -50 1006 -30
rect 1024 -44 1026 -30
rect 1034 -44 1036 -30
rect 1075 -36 1077 -30
rect 1085 -36 1087 -30
rect 1044 -47 1046 -37
rect 1054 -50 1056 -37
rect 1095 -39 1097 -30
rect 1123 -43 1125 -32
rect 1130 -43 1132 -32
rect 1143 -41 1145 -32
rect 1163 -50 1165 -37
rect 1173 -47 1175 -37
rect 1183 -44 1185 -30
rect 1193 -44 1195 -30
rect 1213 -50 1215 -30
rect 1220 -50 1222 -30
rect 1231 -50 1233 -36
rect 1253 -50 1255 -36
rect 1264 -50 1266 -30
rect 1271 -50 1273 -30
rect 1291 -44 1293 -30
rect 1301 -44 1303 -30
rect 1342 -36 1344 -30
rect 1352 -36 1354 -30
rect 1311 -47 1313 -37
rect 1321 -50 1323 -37
rect 1362 -39 1364 -30
rect 1390 -43 1392 -32
rect 1397 -43 1399 -32
rect 1410 -41 1412 -32
rect 1430 -50 1432 -37
rect 1440 -47 1442 -37
rect 1450 -44 1452 -30
rect 1460 -44 1462 -30
rect 1480 -50 1482 -30
rect 1487 -50 1489 -30
rect 1498 -50 1500 -36
rect 1520 -50 1522 -36
rect 1531 -50 1533 -30
rect 1538 -50 1540 -30
rect 1558 -44 1560 -30
rect 1568 -44 1570 -30
rect 1609 -36 1611 -30
rect 1619 -36 1621 -30
rect 1578 -47 1580 -37
rect 1588 -50 1590 -37
rect 1629 -39 1631 -30
rect 1657 -43 1659 -32
rect 1664 -43 1666 -32
rect 1677 -41 1679 -32
rect 1697 -50 1699 -37
rect 1707 -47 1709 -37
rect 1717 -44 1719 -30
rect 1727 -44 1729 -30
rect 1747 -50 1749 -30
rect 1754 -50 1756 -30
rect 1765 -50 1767 -36
rect 1787 -50 1789 -36
rect 1798 -50 1800 -30
rect 1805 -50 1807 -30
rect 1825 -44 1827 -30
rect 1835 -44 1837 -30
rect 1876 -36 1878 -30
rect 1886 -36 1888 -30
rect 1845 -47 1847 -37
rect 1855 -50 1857 -37
rect 1896 -39 1898 -30
rect 1919 -39 1921 -30
rect 1935 -44 1937 -35
rect 1945 -44 1947 -35
rect 1955 -47 1957 -35
rect 1962 -47 1964 -35
rect 1983 -50 1985 -37
rect 1993 -47 1995 -37
rect 2003 -44 2005 -30
rect 2013 -44 2015 -30
rect 2033 -50 2035 -30
rect 2040 -50 2042 -30
rect 2051 -50 2053 -36
rect 2073 -50 2075 -36
rect 2084 -50 2086 -30
rect 2091 -50 2093 -30
rect 2111 -44 2113 -30
rect 2121 -44 2123 -30
rect 2162 -36 2164 -30
rect 2172 -36 2174 -30
rect 2131 -47 2133 -37
rect 2141 -50 2143 -37
rect 2182 -39 2184 -30
rect 2206 -42 2208 -36
rect 2216 -44 2218 -36
rect 2223 -44 2225 -36
rect 2233 -44 2235 -36
rect 2240 -44 2242 -36
rect 2250 -44 2252 -35
rect 2274 -42 2276 -36
rect 2284 -44 2286 -36
rect 2291 -44 2293 -36
rect 2301 -44 2303 -36
rect 2308 -44 2310 -36
rect 2318 -44 2320 -35
rect 15 -80 17 -69
rect 22 -80 24 -69
rect 35 -80 37 -71
rect 55 -80 57 -69
rect 62 -80 64 -69
rect 75 -80 77 -71
rect 95 -75 97 -62
rect 105 -75 107 -65
rect 115 -82 117 -68
rect 125 -82 127 -68
rect 145 -82 147 -62
rect 152 -82 154 -62
rect 163 -76 165 -62
rect 185 -76 187 -62
rect 196 -82 198 -62
rect 203 -82 205 -62
rect 223 -82 225 -68
rect 233 -82 235 -68
rect 243 -75 245 -65
rect 253 -75 255 -62
rect 274 -82 276 -76
rect 284 -82 286 -76
rect 294 -82 296 -73
rect 322 -80 324 -69
rect 329 -80 331 -69
rect 342 -80 344 -71
rect 362 -75 364 -62
rect 372 -75 374 -65
rect 382 -82 384 -68
rect 392 -82 394 -68
rect 412 -82 414 -62
rect 419 -82 421 -62
rect 430 -76 432 -62
rect 452 -76 454 -62
rect 463 -82 465 -62
rect 470 -82 472 -62
rect 490 -82 492 -68
rect 500 -82 502 -68
rect 510 -75 512 -65
rect 520 -75 522 -62
rect 541 -82 543 -76
rect 551 -82 553 -76
rect 561 -82 563 -73
rect 589 -80 591 -69
rect 596 -80 598 -69
rect 609 -80 611 -71
rect 629 -75 631 -62
rect 639 -75 641 -65
rect 649 -82 651 -68
rect 659 -82 661 -68
rect 679 -82 681 -62
rect 686 -82 688 -62
rect 697 -76 699 -62
rect 719 -76 721 -62
rect 730 -82 732 -62
rect 737 -82 739 -62
rect 757 -82 759 -68
rect 767 -82 769 -68
rect 777 -75 779 -65
rect 787 -75 789 -62
rect 808 -82 810 -76
rect 818 -82 820 -76
rect 828 -82 830 -73
rect 856 -80 858 -69
rect 863 -80 865 -69
rect 876 -80 878 -71
rect 896 -75 898 -62
rect 906 -75 908 -65
rect 916 -82 918 -68
rect 926 -82 928 -68
rect 946 -82 948 -62
rect 953 -82 955 -62
rect 964 -76 966 -62
rect 986 -76 988 -62
rect 997 -82 999 -62
rect 1004 -82 1006 -62
rect 1024 -82 1026 -68
rect 1034 -82 1036 -68
rect 1044 -75 1046 -65
rect 1054 -75 1056 -62
rect 1075 -82 1077 -76
rect 1085 -82 1087 -76
rect 1095 -82 1097 -73
rect 1123 -80 1125 -69
rect 1130 -80 1132 -69
rect 1143 -80 1145 -71
rect 1163 -75 1165 -62
rect 1173 -75 1175 -65
rect 1183 -82 1185 -68
rect 1193 -82 1195 -68
rect 1213 -82 1215 -62
rect 1220 -82 1222 -62
rect 1231 -76 1233 -62
rect 1253 -76 1255 -62
rect 1264 -82 1266 -62
rect 1271 -82 1273 -62
rect 1291 -82 1293 -68
rect 1301 -82 1303 -68
rect 1311 -75 1313 -65
rect 1321 -75 1323 -62
rect 1342 -82 1344 -76
rect 1352 -82 1354 -76
rect 1362 -82 1364 -73
rect 1390 -80 1392 -69
rect 1397 -80 1399 -69
rect 1410 -80 1412 -71
rect 1430 -75 1432 -62
rect 1440 -75 1442 -65
rect 1450 -82 1452 -68
rect 1460 -82 1462 -68
rect 1480 -82 1482 -62
rect 1487 -82 1489 -62
rect 1498 -76 1500 -62
rect 1520 -76 1522 -62
rect 1531 -82 1533 -62
rect 1538 -82 1540 -62
rect 1558 -82 1560 -68
rect 1568 -82 1570 -68
rect 1578 -75 1580 -65
rect 1588 -75 1590 -62
rect 1609 -82 1611 -76
rect 1619 -82 1621 -76
rect 1629 -82 1631 -73
rect 1657 -80 1659 -69
rect 1664 -80 1666 -69
rect 1677 -80 1679 -71
rect 1697 -75 1699 -62
rect 1707 -75 1709 -65
rect 1717 -82 1719 -68
rect 1727 -82 1729 -68
rect 1747 -82 1749 -62
rect 1754 -82 1756 -62
rect 1765 -76 1767 -62
rect 1787 -76 1789 -62
rect 1798 -82 1800 -62
rect 1805 -82 1807 -62
rect 1825 -82 1827 -68
rect 1835 -82 1837 -68
rect 1845 -75 1847 -65
rect 1855 -75 1857 -62
rect 1876 -82 1878 -76
rect 1886 -82 1888 -76
rect 1896 -82 1898 -73
rect 1919 -82 1921 -73
rect 1935 -77 1937 -68
rect 1945 -77 1947 -68
rect 1955 -77 1957 -65
rect 1962 -77 1964 -65
rect 1983 -75 1985 -62
rect 1993 -75 1995 -65
rect 2003 -82 2005 -68
rect 2013 -82 2015 -68
rect 2033 -82 2035 -62
rect 2040 -82 2042 -62
rect 2051 -76 2053 -62
rect 2073 -76 2075 -62
rect 2084 -82 2086 -62
rect 2091 -82 2093 -62
rect 2111 -82 2113 -68
rect 2121 -82 2123 -68
rect 2131 -75 2133 -65
rect 2141 -75 2143 -62
rect 2162 -82 2164 -76
rect 2172 -82 2174 -76
rect 2182 -82 2184 -73
rect 2206 -76 2208 -70
rect 2216 -76 2218 -68
rect 2223 -76 2225 -68
rect 2233 -76 2235 -68
rect 2240 -76 2242 -68
rect 2250 -77 2252 -68
rect 2274 -76 2276 -70
rect 2284 -76 2286 -68
rect 2291 -76 2293 -68
rect 2301 -76 2303 -68
rect 2308 -76 2310 -68
rect 2318 -77 2320 -68
rect 15 -187 17 -176
rect 22 -187 24 -176
rect 35 -185 37 -176
rect 55 -187 57 -176
rect 62 -187 64 -176
rect 75 -185 77 -176
rect 95 -194 97 -181
rect 105 -191 107 -181
rect 115 -188 117 -174
rect 125 -188 127 -174
rect 145 -194 147 -174
rect 152 -194 154 -174
rect 163 -194 165 -180
rect 185 -194 187 -180
rect 196 -194 198 -174
rect 203 -194 205 -174
rect 223 -188 225 -174
rect 233 -188 235 -174
rect 274 -180 276 -174
rect 284 -180 286 -174
rect 243 -191 245 -181
rect 253 -194 255 -181
rect 294 -183 296 -174
rect 322 -187 324 -176
rect 329 -187 331 -176
rect 342 -185 344 -176
rect 362 -194 364 -181
rect 372 -191 374 -181
rect 382 -188 384 -174
rect 392 -188 394 -174
rect 412 -194 414 -174
rect 419 -194 421 -174
rect 430 -194 432 -180
rect 452 -194 454 -180
rect 463 -194 465 -174
rect 470 -194 472 -174
rect 490 -188 492 -174
rect 500 -188 502 -174
rect 541 -180 543 -174
rect 551 -180 553 -174
rect 510 -191 512 -181
rect 520 -194 522 -181
rect 561 -183 563 -174
rect 589 -187 591 -176
rect 596 -187 598 -176
rect 609 -185 611 -176
rect 629 -194 631 -181
rect 639 -191 641 -181
rect 649 -188 651 -174
rect 659 -188 661 -174
rect 679 -194 681 -174
rect 686 -194 688 -174
rect 697 -194 699 -180
rect 719 -194 721 -180
rect 730 -194 732 -174
rect 737 -194 739 -174
rect 757 -188 759 -174
rect 767 -188 769 -174
rect 808 -180 810 -174
rect 818 -180 820 -174
rect 777 -191 779 -181
rect 787 -194 789 -181
rect 828 -183 830 -174
rect 856 -187 858 -176
rect 863 -187 865 -176
rect 876 -185 878 -176
rect 896 -194 898 -181
rect 906 -191 908 -181
rect 916 -188 918 -174
rect 926 -188 928 -174
rect 946 -194 948 -174
rect 953 -194 955 -174
rect 964 -194 966 -180
rect 986 -194 988 -180
rect 997 -194 999 -174
rect 1004 -194 1006 -174
rect 1024 -188 1026 -174
rect 1034 -188 1036 -174
rect 1075 -180 1077 -174
rect 1085 -180 1087 -174
rect 1044 -191 1046 -181
rect 1054 -194 1056 -181
rect 1095 -183 1097 -174
rect 1123 -187 1125 -176
rect 1130 -187 1132 -176
rect 1143 -185 1145 -176
rect 1163 -194 1165 -181
rect 1173 -191 1175 -181
rect 1183 -188 1185 -174
rect 1193 -188 1195 -174
rect 1213 -194 1215 -174
rect 1220 -194 1222 -174
rect 1231 -194 1233 -180
rect 1253 -194 1255 -180
rect 1264 -194 1266 -174
rect 1271 -194 1273 -174
rect 1291 -188 1293 -174
rect 1301 -188 1303 -174
rect 1342 -180 1344 -174
rect 1352 -180 1354 -174
rect 1311 -191 1313 -181
rect 1321 -194 1323 -181
rect 1362 -183 1364 -174
rect 1390 -187 1392 -176
rect 1397 -187 1399 -176
rect 1410 -185 1412 -176
rect 1430 -194 1432 -181
rect 1440 -191 1442 -181
rect 1450 -188 1452 -174
rect 1460 -188 1462 -174
rect 1480 -194 1482 -174
rect 1487 -194 1489 -174
rect 1498 -194 1500 -180
rect 1520 -194 1522 -180
rect 1531 -194 1533 -174
rect 1538 -194 1540 -174
rect 1558 -188 1560 -174
rect 1568 -188 1570 -174
rect 1609 -180 1611 -174
rect 1619 -180 1621 -174
rect 1578 -191 1580 -181
rect 1588 -194 1590 -181
rect 1629 -183 1631 -174
rect 1657 -187 1659 -176
rect 1664 -187 1666 -176
rect 1677 -185 1679 -176
rect 1697 -194 1699 -181
rect 1707 -191 1709 -181
rect 1717 -188 1719 -174
rect 1727 -188 1729 -174
rect 1747 -194 1749 -174
rect 1754 -194 1756 -174
rect 1765 -194 1767 -180
rect 1787 -194 1789 -180
rect 1798 -194 1800 -174
rect 1805 -194 1807 -174
rect 1825 -188 1827 -174
rect 1835 -188 1837 -174
rect 1876 -180 1878 -174
rect 1886 -180 1888 -174
rect 1845 -191 1847 -181
rect 1855 -194 1857 -181
rect 1896 -183 1898 -174
rect 1919 -183 1921 -174
rect 1935 -188 1937 -179
rect 1945 -188 1947 -179
rect 1955 -191 1957 -179
rect 1962 -191 1964 -179
rect 1983 -194 1985 -181
rect 1993 -191 1995 -181
rect 2003 -188 2005 -174
rect 2013 -188 2015 -174
rect 2033 -194 2035 -174
rect 2040 -194 2042 -174
rect 2051 -194 2053 -180
rect 2073 -194 2075 -180
rect 2084 -194 2086 -174
rect 2091 -194 2093 -174
rect 2111 -188 2113 -174
rect 2121 -188 2123 -174
rect 2162 -180 2164 -174
rect 2172 -180 2174 -174
rect 2131 -191 2133 -181
rect 2141 -194 2143 -181
rect 2182 -183 2184 -174
rect 2206 -186 2208 -180
rect 2216 -188 2218 -180
rect 2223 -188 2225 -180
rect 2233 -188 2235 -180
rect 2240 -188 2242 -180
rect 2250 -188 2252 -179
rect 2274 -186 2276 -180
rect 2284 -188 2286 -180
rect 2291 -188 2293 -180
rect 2301 -188 2303 -180
rect 2308 -188 2310 -180
rect 2318 -188 2320 -179
rect 15 -224 17 -213
rect 22 -224 24 -213
rect 35 -224 37 -215
rect 55 -224 57 -213
rect 62 -224 64 -213
rect 75 -224 77 -215
rect 95 -219 97 -206
rect 105 -219 107 -209
rect 115 -226 117 -212
rect 125 -226 127 -212
rect 145 -226 147 -206
rect 152 -226 154 -206
rect 163 -220 165 -206
rect 185 -220 187 -206
rect 196 -226 198 -206
rect 203 -226 205 -206
rect 223 -226 225 -212
rect 233 -226 235 -212
rect 243 -219 245 -209
rect 253 -219 255 -206
rect 274 -226 276 -220
rect 284 -226 286 -220
rect 294 -226 296 -217
rect 322 -224 324 -213
rect 329 -224 331 -213
rect 342 -224 344 -215
rect 362 -219 364 -206
rect 372 -219 374 -209
rect 382 -226 384 -212
rect 392 -226 394 -212
rect 412 -226 414 -206
rect 419 -226 421 -206
rect 430 -220 432 -206
rect 452 -220 454 -206
rect 463 -226 465 -206
rect 470 -226 472 -206
rect 490 -226 492 -212
rect 500 -226 502 -212
rect 510 -219 512 -209
rect 520 -219 522 -206
rect 541 -226 543 -220
rect 551 -226 553 -220
rect 561 -226 563 -217
rect 589 -224 591 -213
rect 596 -224 598 -213
rect 609 -224 611 -215
rect 629 -219 631 -206
rect 639 -219 641 -209
rect 649 -226 651 -212
rect 659 -226 661 -212
rect 679 -226 681 -206
rect 686 -226 688 -206
rect 697 -220 699 -206
rect 719 -220 721 -206
rect 730 -226 732 -206
rect 737 -226 739 -206
rect 757 -226 759 -212
rect 767 -226 769 -212
rect 777 -219 779 -209
rect 787 -219 789 -206
rect 808 -226 810 -220
rect 818 -226 820 -220
rect 828 -226 830 -217
rect 856 -224 858 -213
rect 863 -224 865 -213
rect 876 -224 878 -215
rect 896 -219 898 -206
rect 906 -219 908 -209
rect 916 -226 918 -212
rect 926 -226 928 -212
rect 946 -226 948 -206
rect 953 -226 955 -206
rect 964 -220 966 -206
rect 986 -220 988 -206
rect 997 -226 999 -206
rect 1004 -226 1006 -206
rect 1024 -226 1026 -212
rect 1034 -226 1036 -212
rect 1044 -219 1046 -209
rect 1054 -219 1056 -206
rect 1075 -226 1077 -220
rect 1085 -226 1087 -220
rect 1095 -226 1097 -217
rect 1123 -224 1125 -213
rect 1130 -224 1132 -213
rect 1143 -224 1145 -215
rect 1163 -219 1165 -206
rect 1173 -219 1175 -209
rect 1183 -226 1185 -212
rect 1193 -226 1195 -212
rect 1213 -226 1215 -206
rect 1220 -226 1222 -206
rect 1231 -220 1233 -206
rect 1253 -220 1255 -206
rect 1264 -226 1266 -206
rect 1271 -226 1273 -206
rect 1291 -226 1293 -212
rect 1301 -226 1303 -212
rect 1311 -219 1313 -209
rect 1321 -219 1323 -206
rect 1342 -226 1344 -220
rect 1352 -226 1354 -220
rect 1362 -226 1364 -217
rect 1390 -224 1392 -213
rect 1397 -224 1399 -213
rect 1410 -224 1412 -215
rect 1430 -219 1432 -206
rect 1440 -219 1442 -209
rect 1450 -226 1452 -212
rect 1460 -226 1462 -212
rect 1480 -226 1482 -206
rect 1487 -226 1489 -206
rect 1498 -220 1500 -206
rect 1520 -220 1522 -206
rect 1531 -226 1533 -206
rect 1538 -226 1540 -206
rect 1558 -226 1560 -212
rect 1568 -226 1570 -212
rect 1578 -219 1580 -209
rect 1588 -219 1590 -206
rect 1609 -226 1611 -220
rect 1619 -226 1621 -220
rect 1629 -226 1631 -217
rect 1657 -224 1659 -213
rect 1664 -224 1666 -213
rect 1677 -224 1679 -215
rect 1697 -219 1699 -206
rect 1707 -219 1709 -209
rect 1717 -226 1719 -212
rect 1727 -226 1729 -212
rect 1747 -226 1749 -206
rect 1754 -226 1756 -206
rect 1765 -220 1767 -206
rect 1787 -220 1789 -206
rect 1798 -226 1800 -206
rect 1805 -226 1807 -206
rect 1825 -226 1827 -212
rect 1835 -226 1837 -212
rect 1845 -219 1847 -209
rect 1855 -219 1857 -206
rect 1876 -226 1878 -220
rect 1886 -226 1888 -220
rect 1896 -226 1898 -217
rect 1919 -226 1921 -217
rect 1935 -221 1937 -212
rect 1945 -221 1947 -212
rect 1955 -221 1957 -209
rect 1962 -221 1964 -209
rect 1983 -219 1985 -206
rect 1993 -219 1995 -209
rect 2003 -226 2005 -212
rect 2013 -226 2015 -212
rect 2033 -226 2035 -206
rect 2040 -226 2042 -206
rect 2051 -220 2053 -206
rect 2073 -220 2075 -206
rect 2084 -226 2086 -206
rect 2091 -226 2093 -206
rect 2111 -226 2113 -212
rect 2121 -226 2123 -212
rect 2131 -219 2133 -209
rect 2141 -219 2143 -206
rect 2162 -226 2164 -220
rect 2172 -226 2174 -220
rect 2182 -226 2184 -217
rect 2206 -220 2208 -214
rect 2216 -220 2218 -212
rect 2223 -220 2225 -212
rect 2233 -220 2235 -212
rect 2240 -220 2242 -212
rect 2250 -221 2252 -212
rect 2274 -220 2276 -214
rect 2284 -220 2286 -212
rect 2291 -220 2293 -212
rect 2301 -220 2303 -212
rect 2308 -220 2310 -212
rect 2318 -221 2320 -212
<< pmos >>
rect 15 278 17 291
rect 25 278 27 291
rect 35 271 37 289
rect 55 278 57 291
rect 65 278 67 291
rect 75 271 77 289
rect 95 273 97 298
rect 108 273 110 286
rect 118 270 120 295
rect 125 270 127 295
rect 143 270 145 298
rect 153 270 155 298
rect 163 270 165 298
rect 185 270 187 298
rect 195 270 197 298
rect 205 270 207 298
rect 223 270 225 295
rect 230 270 232 295
rect 240 273 242 286
rect 253 273 255 298
rect 274 277 276 298
rect 281 277 283 298
rect 294 270 296 288
rect 322 278 324 291
rect 332 278 334 291
rect 342 271 344 289
rect 362 273 364 298
rect 375 273 377 286
rect 385 270 387 295
rect 392 270 394 295
rect 410 270 412 298
rect 420 270 422 298
rect 430 270 432 298
rect 452 270 454 298
rect 462 270 464 298
rect 472 270 474 298
rect 490 270 492 295
rect 497 270 499 295
rect 507 273 509 286
rect 520 273 522 298
rect 541 277 543 298
rect 548 277 550 298
rect 561 270 563 288
rect 589 278 591 291
rect 599 278 601 291
rect 609 271 611 289
rect 629 273 631 298
rect 642 273 644 286
rect 652 270 654 295
rect 659 270 661 295
rect 677 270 679 298
rect 687 270 689 298
rect 697 270 699 298
rect 719 270 721 298
rect 729 270 731 298
rect 739 270 741 298
rect 757 270 759 295
rect 764 270 766 295
rect 774 273 776 286
rect 787 273 789 298
rect 808 277 810 298
rect 815 277 817 298
rect 828 270 830 288
rect 856 278 858 291
rect 866 278 868 291
rect 876 271 878 289
rect 896 273 898 298
rect 909 273 911 286
rect 919 270 921 295
rect 926 270 928 295
rect 944 270 946 298
rect 954 270 956 298
rect 964 270 966 298
rect 986 270 988 298
rect 996 270 998 298
rect 1006 270 1008 298
rect 1024 270 1026 295
rect 1031 270 1033 295
rect 1041 273 1043 286
rect 1054 273 1056 298
rect 1075 277 1077 298
rect 1082 277 1084 298
rect 1095 270 1097 288
rect 1123 278 1125 291
rect 1133 278 1135 291
rect 1143 271 1145 289
rect 1163 273 1165 298
rect 1176 273 1178 286
rect 1186 270 1188 295
rect 1193 270 1195 295
rect 1211 270 1213 298
rect 1221 270 1223 298
rect 1231 270 1233 298
rect 1253 270 1255 298
rect 1263 270 1265 298
rect 1273 270 1275 298
rect 1291 270 1293 295
rect 1298 270 1300 295
rect 1308 273 1310 286
rect 1321 273 1323 298
rect 1342 277 1344 298
rect 1349 277 1351 298
rect 1362 270 1364 288
rect 1390 278 1392 291
rect 1400 278 1402 291
rect 1410 271 1412 289
rect 1430 273 1432 298
rect 1443 273 1445 286
rect 1453 270 1455 295
rect 1460 270 1462 295
rect 1478 270 1480 298
rect 1488 270 1490 298
rect 1498 270 1500 298
rect 1520 270 1522 298
rect 1530 270 1532 298
rect 1540 270 1542 298
rect 1558 270 1560 295
rect 1565 270 1567 295
rect 1575 273 1577 286
rect 1588 273 1590 298
rect 1609 277 1611 298
rect 1616 277 1618 298
rect 1629 270 1631 288
rect 1657 278 1659 291
rect 1667 278 1669 291
rect 1677 271 1679 289
rect 1697 273 1699 298
rect 1710 273 1712 286
rect 1720 270 1722 295
rect 1727 270 1729 295
rect 1745 270 1747 298
rect 1755 270 1757 298
rect 1765 270 1767 298
rect 1787 270 1789 298
rect 1797 270 1799 298
rect 1807 270 1809 298
rect 1825 270 1827 295
rect 1832 270 1834 295
rect 1842 273 1844 286
rect 1855 273 1857 298
rect 1876 277 1878 298
rect 1883 277 1885 298
rect 1896 270 1898 288
rect 1927 271 1929 298
rect 1943 271 1945 289
rect 1953 271 1955 289
rect 1963 271 1965 298
rect 1983 273 1985 298
rect 1996 273 1998 286
rect 2006 270 2008 295
rect 2013 270 2015 295
rect 2031 270 2033 298
rect 2041 270 2043 298
rect 2051 270 2053 298
rect 2073 270 2075 298
rect 2083 270 2085 298
rect 2093 270 2095 298
rect 2111 270 2113 295
rect 2118 270 2120 295
rect 2128 273 2130 286
rect 2141 273 2143 298
rect 2162 277 2164 298
rect 2169 277 2171 298
rect 2182 270 2184 288
rect 2216 282 2218 298
rect 2223 282 2225 298
rect 2233 282 2235 298
rect 2240 282 2242 298
rect 2206 270 2208 278
rect 2250 280 2252 298
rect 2284 282 2286 298
rect 2291 282 2293 298
rect 2301 282 2303 298
rect 2308 282 2310 298
rect 2274 270 2276 278
rect 2318 280 2320 298
rect 15 173 17 186
rect 25 173 27 186
rect 35 175 37 193
rect 55 173 57 186
rect 65 173 67 186
rect 75 175 77 193
rect 95 166 97 191
rect 108 178 110 191
rect 118 169 120 194
rect 125 169 127 194
rect 143 166 145 194
rect 153 166 155 194
rect 163 166 165 194
rect 185 166 187 194
rect 195 166 197 194
rect 205 166 207 194
rect 223 169 225 194
rect 230 169 232 194
rect 240 178 242 191
rect 253 166 255 191
rect 274 166 276 187
rect 281 166 283 187
rect 294 176 296 194
rect 322 173 324 186
rect 332 173 334 186
rect 342 175 344 193
rect 362 166 364 191
rect 375 178 377 191
rect 385 169 387 194
rect 392 169 394 194
rect 410 166 412 194
rect 420 166 422 194
rect 430 166 432 194
rect 452 166 454 194
rect 462 166 464 194
rect 472 166 474 194
rect 490 169 492 194
rect 497 169 499 194
rect 507 178 509 191
rect 520 166 522 191
rect 541 166 543 187
rect 548 166 550 187
rect 561 176 563 194
rect 589 173 591 186
rect 599 173 601 186
rect 609 175 611 193
rect 629 166 631 191
rect 642 178 644 191
rect 652 169 654 194
rect 659 169 661 194
rect 677 166 679 194
rect 687 166 689 194
rect 697 166 699 194
rect 719 166 721 194
rect 729 166 731 194
rect 739 166 741 194
rect 757 169 759 194
rect 764 169 766 194
rect 774 178 776 191
rect 787 166 789 191
rect 808 166 810 187
rect 815 166 817 187
rect 828 176 830 194
rect 856 173 858 186
rect 866 173 868 186
rect 876 175 878 193
rect 896 166 898 191
rect 909 178 911 191
rect 919 169 921 194
rect 926 169 928 194
rect 944 166 946 194
rect 954 166 956 194
rect 964 166 966 194
rect 986 166 988 194
rect 996 166 998 194
rect 1006 166 1008 194
rect 1024 169 1026 194
rect 1031 169 1033 194
rect 1041 178 1043 191
rect 1054 166 1056 191
rect 1075 166 1077 187
rect 1082 166 1084 187
rect 1095 176 1097 194
rect 1123 173 1125 186
rect 1133 173 1135 186
rect 1143 175 1145 193
rect 1163 166 1165 191
rect 1176 178 1178 191
rect 1186 169 1188 194
rect 1193 169 1195 194
rect 1211 166 1213 194
rect 1221 166 1223 194
rect 1231 166 1233 194
rect 1253 166 1255 194
rect 1263 166 1265 194
rect 1273 166 1275 194
rect 1291 169 1293 194
rect 1298 169 1300 194
rect 1308 178 1310 191
rect 1321 166 1323 191
rect 1342 166 1344 187
rect 1349 166 1351 187
rect 1362 176 1364 194
rect 1390 173 1392 186
rect 1400 173 1402 186
rect 1410 175 1412 193
rect 1430 166 1432 191
rect 1443 178 1445 191
rect 1453 169 1455 194
rect 1460 169 1462 194
rect 1478 166 1480 194
rect 1488 166 1490 194
rect 1498 166 1500 194
rect 1520 166 1522 194
rect 1530 166 1532 194
rect 1540 166 1542 194
rect 1558 169 1560 194
rect 1565 169 1567 194
rect 1575 178 1577 191
rect 1588 166 1590 191
rect 1609 166 1611 187
rect 1616 166 1618 187
rect 1629 176 1631 194
rect 1657 173 1659 186
rect 1667 173 1669 186
rect 1677 175 1679 193
rect 1697 166 1699 191
rect 1710 178 1712 191
rect 1720 169 1722 194
rect 1727 169 1729 194
rect 1745 166 1747 194
rect 1755 166 1757 194
rect 1765 166 1767 194
rect 1787 166 1789 194
rect 1797 166 1799 194
rect 1807 166 1809 194
rect 1825 169 1827 194
rect 1832 169 1834 194
rect 1842 178 1844 191
rect 1855 166 1857 191
rect 1876 166 1878 187
rect 1883 166 1885 187
rect 1896 176 1898 194
rect 1927 166 1929 193
rect 1943 175 1945 193
rect 1953 175 1955 193
rect 1963 166 1965 193
rect 1983 166 1985 191
rect 1996 178 1998 191
rect 2006 169 2008 194
rect 2013 169 2015 194
rect 2031 166 2033 194
rect 2041 166 2043 194
rect 2051 166 2053 194
rect 2073 166 2075 194
rect 2083 166 2085 194
rect 2093 166 2095 194
rect 2111 169 2113 194
rect 2118 169 2120 194
rect 2128 178 2130 191
rect 2141 166 2143 191
rect 2162 166 2164 187
rect 2169 166 2171 187
rect 2182 176 2184 194
rect 2206 186 2208 194
rect 2274 186 2276 194
rect 2216 166 2218 182
rect 2223 166 2225 182
rect 2233 166 2235 182
rect 2240 166 2242 182
rect 2250 166 2252 184
rect 2284 166 2286 182
rect 2291 166 2293 182
rect 2301 166 2303 182
rect 2308 166 2310 182
rect 2318 166 2320 184
rect 15 134 17 147
rect 25 134 27 147
rect 35 127 37 145
rect 55 134 57 147
rect 65 134 67 147
rect 75 127 77 145
rect 95 129 97 154
rect 108 129 110 142
rect 118 126 120 151
rect 125 126 127 151
rect 143 126 145 154
rect 153 126 155 154
rect 163 126 165 154
rect 185 126 187 154
rect 195 126 197 154
rect 205 126 207 154
rect 223 126 225 151
rect 230 126 232 151
rect 240 129 242 142
rect 253 129 255 154
rect 274 133 276 154
rect 281 133 283 154
rect 294 126 296 144
rect 322 134 324 147
rect 332 134 334 147
rect 342 127 344 145
rect 362 129 364 154
rect 375 129 377 142
rect 385 126 387 151
rect 392 126 394 151
rect 410 126 412 154
rect 420 126 422 154
rect 430 126 432 154
rect 452 126 454 154
rect 462 126 464 154
rect 472 126 474 154
rect 490 126 492 151
rect 497 126 499 151
rect 507 129 509 142
rect 520 129 522 154
rect 541 133 543 154
rect 548 133 550 154
rect 561 126 563 144
rect 589 134 591 147
rect 599 134 601 147
rect 609 127 611 145
rect 629 129 631 154
rect 642 129 644 142
rect 652 126 654 151
rect 659 126 661 151
rect 677 126 679 154
rect 687 126 689 154
rect 697 126 699 154
rect 719 126 721 154
rect 729 126 731 154
rect 739 126 741 154
rect 757 126 759 151
rect 764 126 766 151
rect 774 129 776 142
rect 787 129 789 154
rect 808 133 810 154
rect 815 133 817 154
rect 828 126 830 144
rect 856 134 858 147
rect 866 134 868 147
rect 876 127 878 145
rect 896 129 898 154
rect 909 129 911 142
rect 919 126 921 151
rect 926 126 928 151
rect 944 126 946 154
rect 954 126 956 154
rect 964 126 966 154
rect 986 126 988 154
rect 996 126 998 154
rect 1006 126 1008 154
rect 1024 126 1026 151
rect 1031 126 1033 151
rect 1041 129 1043 142
rect 1054 129 1056 154
rect 1075 133 1077 154
rect 1082 133 1084 154
rect 1095 126 1097 144
rect 1123 134 1125 147
rect 1133 134 1135 147
rect 1143 127 1145 145
rect 1163 129 1165 154
rect 1176 129 1178 142
rect 1186 126 1188 151
rect 1193 126 1195 151
rect 1211 126 1213 154
rect 1221 126 1223 154
rect 1231 126 1233 154
rect 1253 126 1255 154
rect 1263 126 1265 154
rect 1273 126 1275 154
rect 1291 126 1293 151
rect 1298 126 1300 151
rect 1308 129 1310 142
rect 1321 129 1323 154
rect 1342 133 1344 154
rect 1349 133 1351 154
rect 1362 126 1364 144
rect 1390 134 1392 147
rect 1400 134 1402 147
rect 1410 127 1412 145
rect 1430 129 1432 154
rect 1443 129 1445 142
rect 1453 126 1455 151
rect 1460 126 1462 151
rect 1478 126 1480 154
rect 1488 126 1490 154
rect 1498 126 1500 154
rect 1520 126 1522 154
rect 1530 126 1532 154
rect 1540 126 1542 154
rect 1558 126 1560 151
rect 1565 126 1567 151
rect 1575 129 1577 142
rect 1588 129 1590 154
rect 1609 133 1611 154
rect 1616 133 1618 154
rect 1629 126 1631 144
rect 1657 134 1659 147
rect 1667 134 1669 147
rect 1677 127 1679 145
rect 1697 129 1699 154
rect 1710 129 1712 142
rect 1720 126 1722 151
rect 1727 126 1729 151
rect 1745 126 1747 154
rect 1755 126 1757 154
rect 1765 126 1767 154
rect 1787 126 1789 154
rect 1797 126 1799 154
rect 1807 126 1809 154
rect 1825 126 1827 151
rect 1832 126 1834 151
rect 1842 129 1844 142
rect 1855 129 1857 154
rect 1876 133 1878 154
rect 1883 133 1885 154
rect 1896 126 1898 144
rect 1927 127 1929 154
rect 1943 127 1945 145
rect 1953 127 1955 145
rect 1963 127 1965 154
rect 1983 129 1985 154
rect 1996 129 1998 142
rect 2006 126 2008 151
rect 2013 126 2015 151
rect 2031 126 2033 154
rect 2041 126 2043 154
rect 2051 126 2053 154
rect 2073 126 2075 154
rect 2083 126 2085 154
rect 2093 126 2095 154
rect 2111 126 2113 151
rect 2118 126 2120 151
rect 2128 129 2130 142
rect 2141 129 2143 154
rect 2162 133 2164 154
rect 2169 133 2171 154
rect 2182 126 2184 144
rect 2216 138 2218 154
rect 2223 138 2225 154
rect 2233 138 2235 154
rect 2240 138 2242 154
rect 2206 126 2208 134
rect 2250 136 2252 154
rect 2284 138 2286 154
rect 2291 138 2293 154
rect 2301 138 2303 154
rect 2308 138 2310 154
rect 2274 126 2276 134
rect 2318 136 2320 154
rect 15 29 17 42
rect 25 29 27 42
rect 35 31 37 49
rect 55 29 57 42
rect 65 29 67 42
rect 75 31 77 49
rect 95 22 97 47
rect 108 34 110 47
rect 118 25 120 50
rect 125 25 127 50
rect 143 22 145 50
rect 153 22 155 50
rect 163 22 165 50
rect 185 22 187 50
rect 195 22 197 50
rect 205 22 207 50
rect 223 25 225 50
rect 230 25 232 50
rect 240 34 242 47
rect 253 22 255 47
rect 274 22 276 43
rect 281 22 283 43
rect 294 32 296 50
rect 322 29 324 42
rect 332 29 334 42
rect 342 31 344 49
rect 362 22 364 47
rect 375 34 377 47
rect 385 25 387 50
rect 392 25 394 50
rect 410 22 412 50
rect 420 22 422 50
rect 430 22 432 50
rect 452 22 454 50
rect 462 22 464 50
rect 472 22 474 50
rect 490 25 492 50
rect 497 25 499 50
rect 507 34 509 47
rect 520 22 522 47
rect 541 22 543 43
rect 548 22 550 43
rect 561 32 563 50
rect 589 29 591 42
rect 599 29 601 42
rect 609 31 611 49
rect 629 22 631 47
rect 642 34 644 47
rect 652 25 654 50
rect 659 25 661 50
rect 677 22 679 50
rect 687 22 689 50
rect 697 22 699 50
rect 719 22 721 50
rect 729 22 731 50
rect 739 22 741 50
rect 757 25 759 50
rect 764 25 766 50
rect 774 34 776 47
rect 787 22 789 47
rect 808 22 810 43
rect 815 22 817 43
rect 828 32 830 50
rect 856 29 858 42
rect 866 29 868 42
rect 876 31 878 49
rect 896 22 898 47
rect 909 34 911 47
rect 919 25 921 50
rect 926 25 928 50
rect 944 22 946 50
rect 954 22 956 50
rect 964 22 966 50
rect 986 22 988 50
rect 996 22 998 50
rect 1006 22 1008 50
rect 1024 25 1026 50
rect 1031 25 1033 50
rect 1041 34 1043 47
rect 1054 22 1056 47
rect 1075 22 1077 43
rect 1082 22 1084 43
rect 1095 32 1097 50
rect 1123 29 1125 42
rect 1133 29 1135 42
rect 1143 31 1145 49
rect 1163 22 1165 47
rect 1176 34 1178 47
rect 1186 25 1188 50
rect 1193 25 1195 50
rect 1211 22 1213 50
rect 1221 22 1223 50
rect 1231 22 1233 50
rect 1253 22 1255 50
rect 1263 22 1265 50
rect 1273 22 1275 50
rect 1291 25 1293 50
rect 1298 25 1300 50
rect 1308 34 1310 47
rect 1321 22 1323 47
rect 1342 22 1344 43
rect 1349 22 1351 43
rect 1362 32 1364 50
rect 1390 29 1392 42
rect 1400 29 1402 42
rect 1410 31 1412 49
rect 1430 22 1432 47
rect 1443 34 1445 47
rect 1453 25 1455 50
rect 1460 25 1462 50
rect 1478 22 1480 50
rect 1488 22 1490 50
rect 1498 22 1500 50
rect 1520 22 1522 50
rect 1530 22 1532 50
rect 1540 22 1542 50
rect 1558 25 1560 50
rect 1565 25 1567 50
rect 1575 34 1577 47
rect 1588 22 1590 47
rect 1609 22 1611 43
rect 1616 22 1618 43
rect 1629 32 1631 50
rect 1657 29 1659 42
rect 1667 29 1669 42
rect 1677 31 1679 49
rect 1697 22 1699 47
rect 1710 34 1712 47
rect 1720 25 1722 50
rect 1727 25 1729 50
rect 1745 22 1747 50
rect 1755 22 1757 50
rect 1765 22 1767 50
rect 1787 22 1789 50
rect 1797 22 1799 50
rect 1807 22 1809 50
rect 1825 25 1827 50
rect 1832 25 1834 50
rect 1842 34 1844 47
rect 1855 22 1857 47
rect 1876 22 1878 43
rect 1883 22 1885 43
rect 1896 32 1898 50
rect 1927 22 1929 49
rect 1943 31 1945 49
rect 1953 31 1955 49
rect 1963 22 1965 49
rect 1983 22 1985 47
rect 1996 34 1998 47
rect 2006 25 2008 50
rect 2013 25 2015 50
rect 2031 22 2033 50
rect 2041 22 2043 50
rect 2051 22 2053 50
rect 2073 22 2075 50
rect 2083 22 2085 50
rect 2093 22 2095 50
rect 2111 25 2113 50
rect 2118 25 2120 50
rect 2128 34 2130 47
rect 2141 22 2143 47
rect 2162 22 2164 43
rect 2169 22 2171 43
rect 2182 32 2184 50
rect 2206 42 2208 50
rect 2274 42 2276 50
rect 2216 22 2218 38
rect 2223 22 2225 38
rect 2233 22 2235 38
rect 2240 22 2242 38
rect 2250 22 2252 40
rect 2284 22 2286 38
rect 2291 22 2293 38
rect 2301 22 2303 38
rect 2308 22 2310 38
rect 2318 22 2320 40
rect 15 -10 17 3
rect 25 -10 27 3
rect 35 -17 37 1
rect 55 -10 57 3
rect 65 -10 67 3
rect 75 -17 77 1
rect 95 -15 97 10
rect 108 -15 110 -2
rect 118 -18 120 7
rect 125 -18 127 7
rect 143 -18 145 10
rect 153 -18 155 10
rect 163 -18 165 10
rect 185 -18 187 10
rect 195 -18 197 10
rect 205 -18 207 10
rect 223 -18 225 7
rect 230 -18 232 7
rect 240 -15 242 -2
rect 253 -15 255 10
rect 274 -11 276 10
rect 281 -11 283 10
rect 294 -18 296 0
rect 322 -10 324 3
rect 332 -10 334 3
rect 342 -17 344 1
rect 362 -15 364 10
rect 375 -15 377 -2
rect 385 -18 387 7
rect 392 -18 394 7
rect 410 -18 412 10
rect 420 -18 422 10
rect 430 -18 432 10
rect 452 -18 454 10
rect 462 -18 464 10
rect 472 -18 474 10
rect 490 -18 492 7
rect 497 -18 499 7
rect 507 -15 509 -2
rect 520 -15 522 10
rect 541 -11 543 10
rect 548 -11 550 10
rect 561 -18 563 0
rect 589 -10 591 3
rect 599 -10 601 3
rect 609 -17 611 1
rect 629 -15 631 10
rect 642 -15 644 -2
rect 652 -18 654 7
rect 659 -18 661 7
rect 677 -18 679 10
rect 687 -18 689 10
rect 697 -18 699 10
rect 719 -18 721 10
rect 729 -18 731 10
rect 739 -18 741 10
rect 757 -18 759 7
rect 764 -18 766 7
rect 774 -15 776 -2
rect 787 -15 789 10
rect 808 -11 810 10
rect 815 -11 817 10
rect 828 -18 830 0
rect 856 -10 858 3
rect 866 -10 868 3
rect 876 -17 878 1
rect 896 -15 898 10
rect 909 -15 911 -2
rect 919 -18 921 7
rect 926 -18 928 7
rect 944 -18 946 10
rect 954 -18 956 10
rect 964 -18 966 10
rect 986 -18 988 10
rect 996 -18 998 10
rect 1006 -18 1008 10
rect 1024 -18 1026 7
rect 1031 -18 1033 7
rect 1041 -15 1043 -2
rect 1054 -15 1056 10
rect 1075 -11 1077 10
rect 1082 -11 1084 10
rect 1095 -18 1097 0
rect 1123 -10 1125 3
rect 1133 -10 1135 3
rect 1143 -17 1145 1
rect 1163 -15 1165 10
rect 1176 -15 1178 -2
rect 1186 -18 1188 7
rect 1193 -18 1195 7
rect 1211 -18 1213 10
rect 1221 -18 1223 10
rect 1231 -18 1233 10
rect 1253 -18 1255 10
rect 1263 -18 1265 10
rect 1273 -18 1275 10
rect 1291 -18 1293 7
rect 1298 -18 1300 7
rect 1308 -15 1310 -2
rect 1321 -15 1323 10
rect 1342 -11 1344 10
rect 1349 -11 1351 10
rect 1362 -18 1364 0
rect 1390 -10 1392 3
rect 1400 -10 1402 3
rect 1410 -17 1412 1
rect 1430 -15 1432 10
rect 1443 -15 1445 -2
rect 1453 -18 1455 7
rect 1460 -18 1462 7
rect 1478 -18 1480 10
rect 1488 -18 1490 10
rect 1498 -18 1500 10
rect 1520 -18 1522 10
rect 1530 -18 1532 10
rect 1540 -18 1542 10
rect 1558 -18 1560 7
rect 1565 -18 1567 7
rect 1575 -15 1577 -2
rect 1588 -15 1590 10
rect 1609 -11 1611 10
rect 1616 -11 1618 10
rect 1629 -18 1631 0
rect 1657 -10 1659 3
rect 1667 -10 1669 3
rect 1677 -17 1679 1
rect 1697 -15 1699 10
rect 1710 -15 1712 -2
rect 1720 -18 1722 7
rect 1727 -18 1729 7
rect 1745 -18 1747 10
rect 1755 -18 1757 10
rect 1765 -18 1767 10
rect 1787 -18 1789 10
rect 1797 -18 1799 10
rect 1807 -18 1809 10
rect 1825 -18 1827 7
rect 1832 -18 1834 7
rect 1842 -15 1844 -2
rect 1855 -15 1857 10
rect 1876 -11 1878 10
rect 1883 -11 1885 10
rect 1896 -18 1898 0
rect 1927 -17 1929 10
rect 1943 -17 1945 1
rect 1953 -17 1955 1
rect 1963 -17 1965 10
rect 1983 -15 1985 10
rect 1996 -15 1998 -2
rect 2006 -18 2008 7
rect 2013 -18 2015 7
rect 2031 -18 2033 10
rect 2041 -18 2043 10
rect 2051 -18 2053 10
rect 2073 -18 2075 10
rect 2083 -18 2085 10
rect 2093 -18 2095 10
rect 2111 -18 2113 7
rect 2118 -18 2120 7
rect 2128 -15 2130 -2
rect 2141 -15 2143 10
rect 2162 -11 2164 10
rect 2169 -11 2171 10
rect 2182 -18 2184 0
rect 2216 -6 2218 10
rect 2223 -6 2225 10
rect 2233 -6 2235 10
rect 2240 -6 2242 10
rect 2206 -18 2208 -10
rect 2250 -8 2252 10
rect 2284 -6 2286 10
rect 2291 -6 2293 10
rect 2301 -6 2303 10
rect 2308 -6 2310 10
rect 2274 -18 2276 -10
rect 2318 -8 2320 10
rect 15 -115 17 -102
rect 25 -115 27 -102
rect 35 -113 37 -95
rect 55 -115 57 -102
rect 65 -115 67 -102
rect 75 -113 77 -95
rect 95 -122 97 -97
rect 108 -110 110 -97
rect 118 -119 120 -94
rect 125 -119 127 -94
rect 143 -122 145 -94
rect 153 -122 155 -94
rect 163 -122 165 -94
rect 185 -122 187 -94
rect 195 -122 197 -94
rect 205 -122 207 -94
rect 223 -119 225 -94
rect 230 -119 232 -94
rect 240 -110 242 -97
rect 253 -122 255 -97
rect 274 -122 276 -101
rect 281 -122 283 -101
rect 294 -112 296 -94
rect 322 -115 324 -102
rect 332 -115 334 -102
rect 342 -113 344 -95
rect 362 -122 364 -97
rect 375 -110 377 -97
rect 385 -119 387 -94
rect 392 -119 394 -94
rect 410 -122 412 -94
rect 420 -122 422 -94
rect 430 -122 432 -94
rect 452 -122 454 -94
rect 462 -122 464 -94
rect 472 -122 474 -94
rect 490 -119 492 -94
rect 497 -119 499 -94
rect 507 -110 509 -97
rect 520 -122 522 -97
rect 541 -122 543 -101
rect 548 -122 550 -101
rect 561 -112 563 -94
rect 589 -115 591 -102
rect 599 -115 601 -102
rect 609 -113 611 -95
rect 629 -122 631 -97
rect 642 -110 644 -97
rect 652 -119 654 -94
rect 659 -119 661 -94
rect 677 -122 679 -94
rect 687 -122 689 -94
rect 697 -122 699 -94
rect 719 -122 721 -94
rect 729 -122 731 -94
rect 739 -122 741 -94
rect 757 -119 759 -94
rect 764 -119 766 -94
rect 774 -110 776 -97
rect 787 -122 789 -97
rect 808 -122 810 -101
rect 815 -122 817 -101
rect 828 -112 830 -94
rect 856 -115 858 -102
rect 866 -115 868 -102
rect 876 -113 878 -95
rect 896 -122 898 -97
rect 909 -110 911 -97
rect 919 -119 921 -94
rect 926 -119 928 -94
rect 944 -122 946 -94
rect 954 -122 956 -94
rect 964 -122 966 -94
rect 986 -122 988 -94
rect 996 -122 998 -94
rect 1006 -122 1008 -94
rect 1024 -119 1026 -94
rect 1031 -119 1033 -94
rect 1041 -110 1043 -97
rect 1054 -122 1056 -97
rect 1075 -122 1077 -101
rect 1082 -122 1084 -101
rect 1095 -112 1097 -94
rect 1123 -115 1125 -102
rect 1133 -115 1135 -102
rect 1143 -113 1145 -95
rect 1163 -122 1165 -97
rect 1176 -110 1178 -97
rect 1186 -119 1188 -94
rect 1193 -119 1195 -94
rect 1211 -122 1213 -94
rect 1221 -122 1223 -94
rect 1231 -122 1233 -94
rect 1253 -122 1255 -94
rect 1263 -122 1265 -94
rect 1273 -122 1275 -94
rect 1291 -119 1293 -94
rect 1298 -119 1300 -94
rect 1308 -110 1310 -97
rect 1321 -122 1323 -97
rect 1342 -122 1344 -101
rect 1349 -122 1351 -101
rect 1362 -112 1364 -94
rect 1390 -115 1392 -102
rect 1400 -115 1402 -102
rect 1410 -113 1412 -95
rect 1430 -122 1432 -97
rect 1443 -110 1445 -97
rect 1453 -119 1455 -94
rect 1460 -119 1462 -94
rect 1478 -122 1480 -94
rect 1488 -122 1490 -94
rect 1498 -122 1500 -94
rect 1520 -122 1522 -94
rect 1530 -122 1532 -94
rect 1540 -122 1542 -94
rect 1558 -119 1560 -94
rect 1565 -119 1567 -94
rect 1575 -110 1577 -97
rect 1588 -122 1590 -97
rect 1609 -122 1611 -101
rect 1616 -122 1618 -101
rect 1629 -112 1631 -94
rect 1657 -115 1659 -102
rect 1667 -115 1669 -102
rect 1677 -113 1679 -95
rect 1697 -122 1699 -97
rect 1710 -110 1712 -97
rect 1720 -119 1722 -94
rect 1727 -119 1729 -94
rect 1745 -122 1747 -94
rect 1755 -122 1757 -94
rect 1765 -122 1767 -94
rect 1787 -122 1789 -94
rect 1797 -122 1799 -94
rect 1807 -122 1809 -94
rect 1825 -119 1827 -94
rect 1832 -119 1834 -94
rect 1842 -110 1844 -97
rect 1855 -122 1857 -97
rect 1876 -122 1878 -101
rect 1883 -122 1885 -101
rect 1896 -112 1898 -94
rect 1927 -122 1929 -95
rect 1943 -113 1945 -95
rect 1953 -113 1955 -95
rect 1963 -122 1965 -95
rect 1983 -122 1985 -97
rect 1996 -110 1998 -97
rect 2006 -119 2008 -94
rect 2013 -119 2015 -94
rect 2031 -122 2033 -94
rect 2041 -122 2043 -94
rect 2051 -122 2053 -94
rect 2073 -122 2075 -94
rect 2083 -122 2085 -94
rect 2093 -122 2095 -94
rect 2111 -119 2113 -94
rect 2118 -119 2120 -94
rect 2128 -110 2130 -97
rect 2141 -122 2143 -97
rect 2162 -122 2164 -101
rect 2169 -122 2171 -101
rect 2182 -112 2184 -94
rect 2206 -102 2208 -94
rect 2274 -102 2276 -94
rect 2216 -122 2218 -106
rect 2223 -122 2225 -106
rect 2233 -122 2235 -106
rect 2240 -122 2242 -106
rect 2250 -122 2252 -104
rect 2284 -122 2286 -106
rect 2291 -122 2293 -106
rect 2301 -122 2303 -106
rect 2308 -122 2310 -106
rect 2318 -122 2320 -104
rect 15 -154 17 -141
rect 25 -154 27 -141
rect 35 -161 37 -143
rect 55 -154 57 -141
rect 65 -154 67 -141
rect 75 -161 77 -143
rect 95 -159 97 -134
rect 108 -159 110 -146
rect 118 -162 120 -137
rect 125 -162 127 -137
rect 143 -162 145 -134
rect 153 -162 155 -134
rect 163 -162 165 -134
rect 185 -162 187 -134
rect 195 -162 197 -134
rect 205 -162 207 -134
rect 223 -162 225 -137
rect 230 -162 232 -137
rect 240 -159 242 -146
rect 253 -159 255 -134
rect 274 -155 276 -134
rect 281 -155 283 -134
rect 294 -162 296 -144
rect 322 -154 324 -141
rect 332 -154 334 -141
rect 342 -161 344 -143
rect 362 -159 364 -134
rect 375 -159 377 -146
rect 385 -162 387 -137
rect 392 -162 394 -137
rect 410 -162 412 -134
rect 420 -162 422 -134
rect 430 -162 432 -134
rect 452 -162 454 -134
rect 462 -162 464 -134
rect 472 -162 474 -134
rect 490 -162 492 -137
rect 497 -162 499 -137
rect 507 -159 509 -146
rect 520 -159 522 -134
rect 541 -155 543 -134
rect 548 -155 550 -134
rect 561 -162 563 -144
rect 589 -154 591 -141
rect 599 -154 601 -141
rect 609 -161 611 -143
rect 629 -159 631 -134
rect 642 -159 644 -146
rect 652 -162 654 -137
rect 659 -162 661 -137
rect 677 -162 679 -134
rect 687 -162 689 -134
rect 697 -162 699 -134
rect 719 -162 721 -134
rect 729 -162 731 -134
rect 739 -162 741 -134
rect 757 -162 759 -137
rect 764 -162 766 -137
rect 774 -159 776 -146
rect 787 -159 789 -134
rect 808 -155 810 -134
rect 815 -155 817 -134
rect 828 -162 830 -144
rect 856 -154 858 -141
rect 866 -154 868 -141
rect 876 -161 878 -143
rect 896 -159 898 -134
rect 909 -159 911 -146
rect 919 -162 921 -137
rect 926 -162 928 -137
rect 944 -162 946 -134
rect 954 -162 956 -134
rect 964 -162 966 -134
rect 986 -162 988 -134
rect 996 -162 998 -134
rect 1006 -162 1008 -134
rect 1024 -162 1026 -137
rect 1031 -162 1033 -137
rect 1041 -159 1043 -146
rect 1054 -159 1056 -134
rect 1075 -155 1077 -134
rect 1082 -155 1084 -134
rect 1095 -162 1097 -144
rect 1123 -154 1125 -141
rect 1133 -154 1135 -141
rect 1143 -161 1145 -143
rect 1163 -159 1165 -134
rect 1176 -159 1178 -146
rect 1186 -162 1188 -137
rect 1193 -162 1195 -137
rect 1211 -162 1213 -134
rect 1221 -162 1223 -134
rect 1231 -162 1233 -134
rect 1253 -162 1255 -134
rect 1263 -162 1265 -134
rect 1273 -162 1275 -134
rect 1291 -162 1293 -137
rect 1298 -162 1300 -137
rect 1308 -159 1310 -146
rect 1321 -159 1323 -134
rect 1342 -155 1344 -134
rect 1349 -155 1351 -134
rect 1362 -162 1364 -144
rect 1390 -154 1392 -141
rect 1400 -154 1402 -141
rect 1410 -161 1412 -143
rect 1430 -159 1432 -134
rect 1443 -159 1445 -146
rect 1453 -162 1455 -137
rect 1460 -162 1462 -137
rect 1478 -162 1480 -134
rect 1488 -162 1490 -134
rect 1498 -162 1500 -134
rect 1520 -162 1522 -134
rect 1530 -162 1532 -134
rect 1540 -162 1542 -134
rect 1558 -162 1560 -137
rect 1565 -162 1567 -137
rect 1575 -159 1577 -146
rect 1588 -159 1590 -134
rect 1609 -155 1611 -134
rect 1616 -155 1618 -134
rect 1629 -162 1631 -144
rect 1657 -154 1659 -141
rect 1667 -154 1669 -141
rect 1677 -161 1679 -143
rect 1697 -159 1699 -134
rect 1710 -159 1712 -146
rect 1720 -162 1722 -137
rect 1727 -162 1729 -137
rect 1745 -162 1747 -134
rect 1755 -162 1757 -134
rect 1765 -162 1767 -134
rect 1787 -162 1789 -134
rect 1797 -162 1799 -134
rect 1807 -162 1809 -134
rect 1825 -162 1827 -137
rect 1832 -162 1834 -137
rect 1842 -159 1844 -146
rect 1855 -159 1857 -134
rect 1876 -155 1878 -134
rect 1883 -155 1885 -134
rect 1896 -162 1898 -144
rect 1927 -161 1929 -134
rect 1943 -161 1945 -143
rect 1953 -161 1955 -143
rect 1963 -161 1965 -134
rect 1983 -159 1985 -134
rect 1996 -159 1998 -146
rect 2006 -162 2008 -137
rect 2013 -162 2015 -137
rect 2031 -162 2033 -134
rect 2041 -162 2043 -134
rect 2051 -162 2053 -134
rect 2073 -162 2075 -134
rect 2083 -162 2085 -134
rect 2093 -162 2095 -134
rect 2111 -162 2113 -137
rect 2118 -162 2120 -137
rect 2128 -159 2130 -146
rect 2141 -159 2143 -134
rect 2162 -155 2164 -134
rect 2169 -155 2171 -134
rect 2182 -162 2184 -144
rect 2216 -150 2218 -134
rect 2223 -150 2225 -134
rect 2233 -150 2235 -134
rect 2240 -150 2242 -134
rect 2206 -162 2208 -154
rect 2250 -152 2252 -134
rect 2284 -150 2286 -134
rect 2291 -150 2293 -134
rect 2301 -150 2303 -134
rect 2308 -150 2310 -134
rect 2274 -162 2276 -154
rect 2318 -152 2320 -134
rect 15 -259 17 -246
rect 25 -259 27 -246
rect 35 -257 37 -239
rect 55 -259 57 -246
rect 65 -259 67 -246
rect 75 -257 77 -239
rect 95 -266 97 -241
rect 108 -254 110 -241
rect 118 -263 120 -238
rect 125 -263 127 -238
rect 143 -266 145 -238
rect 153 -266 155 -238
rect 163 -266 165 -238
rect 185 -266 187 -238
rect 195 -266 197 -238
rect 205 -266 207 -238
rect 223 -263 225 -238
rect 230 -263 232 -238
rect 240 -254 242 -241
rect 253 -266 255 -241
rect 274 -266 276 -245
rect 281 -266 283 -245
rect 294 -256 296 -238
rect 322 -259 324 -246
rect 332 -259 334 -246
rect 342 -257 344 -239
rect 362 -266 364 -241
rect 375 -254 377 -241
rect 385 -263 387 -238
rect 392 -263 394 -238
rect 410 -266 412 -238
rect 420 -266 422 -238
rect 430 -266 432 -238
rect 452 -266 454 -238
rect 462 -266 464 -238
rect 472 -266 474 -238
rect 490 -263 492 -238
rect 497 -263 499 -238
rect 507 -254 509 -241
rect 520 -266 522 -241
rect 541 -266 543 -245
rect 548 -266 550 -245
rect 561 -256 563 -238
rect 589 -259 591 -246
rect 599 -259 601 -246
rect 609 -257 611 -239
rect 629 -266 631 -241
rect 642 -254 644 -241
rect 652 -263 654 -238
rect 659 -263 661 -238
rect 677 -266 679 -238
rect 687 -266 689 -238
rect 697 -266 699 -238
rect 719 -266 721 -238
rect 729 -266 731 -238
rect 739 -266 741 -238
rect 757 -263 759 -238
rect 764 -263 766 -238
rect 774 -254 776 -241
rect 787 -266 789 -241
rect 808 -266 810 -245
rect 815 -266 817 -245
rect 828 -256 830 -238
rect 856 -259 858 -246
rect 866 -259 868 -246
rect 876 -257 878 -239
rect 896 -266 898 -241
rect 909 -254 911 -241
rect 919 -263 921 -238
rect 926 -263 928 -238
rect 944 -266 946 -238
rect 954 -266 956 -238
rect 964 -266 966 -238
rect 986 -266 988 -238
rect 996 -266 998 -238
rect 1006 -266 1008 -238
rect 1024 -263 1026 -238
rect 1031 -263 1033 -238
rect 1041 -254 1043 -241
rect 1054 -266 1056 -241
rect 1075 -266 1077 -245
rect 1082 -266 1084 -245
rect 1095 -256 1097 -238
rect 1123 -259 1125 -246
rect 1133 -259 1135 -246
rect 1143 -257 1145 -239
rect 1163 -266 1165 -241
rect 1176 -254 1178 -241
rect 1186 -263 1188 -238
rect 1193 -263 1195 -238
rect 1211 -266 1213 -238
rect 1221 -266 1223 -238
rect 1231 -266 1233 -238
rect 1253 -266 1255 -238
rect 1263 -266 1265 -238
rect 1273 -266 1275 -238
rect 1291 -263 1293 -238
rect 1298 -263 1300 -238
rect 1308 -254 1310 -241
rect 1321 -266 1323 -241
rect 1342 -266 1344 -245
rect 1349 -266 1351 -245
rect 1362 -256 1364 -238
rect 1390 -259 1392 -246
rect 1400 -259 1402 -246
rect 1410 -257 1412 -239
rect 1430 -266 1432 -241
rect 1443 -254 1445 -241
rect 1453 -263 1455 -238
rect 1460 -263 1462 -238
rect 1478 -266 1480 -238
rect 1488 -266 1490 -238
rect 1498 -266 1500 -238
rect 1520 -266 1522 -238
rect 1530 -266 1532 -238
rect 1540 -266 1542 -238
rect 1558 -263 1560 -238
rect 1565 -263 1567 -238
rect 1575 -254 1577 -241
rect 1588 -266 1590 -241
rect 1609 -266 1611 -245
rect 1616 -266 1618 -245
rect 1629 -256 1631 -238
rect 1657 -259 1659 -246
rect 1667 -259 1669 -246
rect 1677 -257 1679 -239
rect 1697 -266 1699 -241
rect 1710 -254 1712 -241
rect 1720 -263 1722 -238
rect 1727 -263 1729 -238
rect 1745 -266 1747 -238
rect 1755 -266 1757 -238
rect 1765 -266 1767 -238
rect 1787 -266 1789 -238
rect 1797 -266 1799 -238
rect 1807 -266 1809 -238
rect 1825 -263 1827 -238
rect 1832 -263 1834 -238
rect 1842 -254 1844 -241
rect 1855 -266 1857 -241
rect 1876 -266 1878 -245
rect 1883 -266 1885 -245
rect 1896 -256 1898 -238
rect 1927 -266 1929 -239
rect 1943 -257 1945 -239
rect 1953 -257 1955 -239
rect 1963 -266 1965 -239
rect 1983 -266 1985 -241
rect 1996 -254 1998 -241
rect 2006 -263 2008 -238
rect 2013 -263 2015 -238
rect 2031 -266 2033 -238
rect 2041 -266 2043 -238
rect 2051 -266 2053 -238
rect 2073 -266 2075 -238
rect 2083 -266 2085 -238
rect 2093 -266 2095 -238
rect 2111 -263 2113 -238
rect 2118 -263 2120 -238
rect 2128 -254 2130 -241
rect 2141 -266 2143 -241
rect 2162 -266 2164 -245
rect 2169 -266 2171 -245
rect 2182 -256 2184 -238
rect 2206 -246 2208 -238
rect 2274 -246 2276 -238
rect 2216 -266 2218 -250
rect 2223 -266 2225 -250
rect 2233 -266 2235 -250
rect 2240 -266 2242 -250
rect 2250 -266 2252 -248
rect 2284 -266 2286 -250
rect 2291 -266 2293 -250
rect 2301 -266 2303 -250
rect 2308 -266 2310 -250
rect 2318 -266 2320 -248
<< polyct0 >>
rect 33 263 35 265
rect 73 263 75 265
rect 103 266 105 268
rect 97 256 99 258
rect 153 263 155 265
rect 163 263 165 265
rect 185 263 187 265
rect 195 263 197 265
rect 245 266 247 268
rect 292 263 294 265
rect 251 256 253 258
rect 340 263 342 265
rect 370 266 372 268
rect 364 256 366 258
rect 420 263 422 265
rect 430 263 432 265
rect 452 263 454 265
rect 462 263 464 265
rect 512 266 514 268
rect 559 263 561 265
rect 518 256 520 258
rect 607 263 609 265
rect 637 266 639 268
rect 631 256 633 258
rect 687 263 689 265
rect 697 263 699 265
rect 719 263 721 265
rect 729 263 731 265
rect 779 266 781 268
rect 826 263 828 265
rect 785 256 787 258
rect 874 263 876 265
rect 904 266 906 268
rect 898 256 900 258
rect 954 263 956 265
rect 964 263 966 265
rect 986 263 988 265
rect 996 263 998 265
rect 1046 266 1048 268
rect 1093 263 1095 265
rect 1052 256 1054 258
rect 1141 263 1143 265
rect 1171 266 1173 268
rect 1165 256 1167 258
rect 1221 263 1223 265
rect 1231 263 1233 265
rect 1253 263 1255 265
rect 1263 263 1265 265
rect 1313 266 1315 268
rect 1360 263 1362 265
rect 1319 256 1321 258
rect 1408 263 1410 265
rect 1438 266 1440 268
rect 1432 256 1434 258
rect 1488 263 1490 265
rect 1498 263 1500 265
rect 1520 263 1522 265
rect 1530 263 1532 265
rect 1580 266 1582 268
rect 1627 263 1629 265
rect 1586 256 1588 258
rect 1675 263 1677 265
rect 1705 266 1707 268
rect 1699 256 1701 258
rect 1755 263 1757 265
rect 1765 263 1767 265
rect 1787 263 1789 265
rect 1797 263 1799 265
rect 1847 266 1849 268
rect 1894 263 1896 265
rect 1951 263 1953 265
rect 1961 264 1963 266
rect 1853 256 1855 258
rect 1991 266 1993 268
rect 1985 256 1987 258
rect 2041 263 2043 265
rect 2051 263 2053 265
rect 2073 263 2075 265
rect 2083 263 2085 265
rect 2133 266 2135 268
rect 2180 263 2182 265
rect 2139 256 2141 258
rect 2224 273 2226 275
rect 2231 257 2233 259
rect 2249 258 2251 260
rect 2292 273 2294 275
rect 2299 257 2301 259
rect 2317 258 2319 260
rect 33 199 35 201
rect 73 199 75 201
rect 97 206 99 208
rect 103 196 105 198
rect 153 199 155 201
rect 163 199 165 201
rect 185 199 187 201
rect 195 199 197 201
rect 251 206 253 208
rect 245 196 247 198
rect 292 199 294 201
rect 340 199 342 201
rect 364 206 366 208
rect 370 196 372 198
rect 420 199 422 201
rect 430 199 432 201
rect 452 199 454 201
rect 462 199 464 201
rect 518 206 520 208
rect 512 196 514 198
rect 559 199 561 201
rect 607 199 609 201
rect 631 206 633 208
rect 637 196 639 198
rect 687 199 689 201
rect 697 199 699 201
rect 719 199 721 201
rect 729 199 731 201
rect 785 206 787 208
rect 779 196 781 198
rect 826 199 828 201
rect 874 199 876 201
rect 898 206 900 208
rect 904 196 906 198
rect 954 199 956 201
rect 964 199 966 201
rect 986 199 988 201
rect 996 199 998 201
rect 1052 206 1054 208
rect 1046 196 1048 198
rect 1093 199 1095 201
rect 1141 199 1143 201
rect 1165 206 1167 208
rect 1171 196 1173 198
rect 1221 199 1223 201
rect 1231 199 1233 201
rect 1253 199 1255 201
rect 1263 199 1265 201
rect 1319 206 1321 208
rect 1313 196 1315 198
rect 1360 199 1362 201
rect 1408 199 1410 201
rect 1432 206 1434 208
rect 1438 196 1440 198
rect 1488 199 1490 201
rect 1498 199 1500 201
rect 1520 199 1522 201
rect 1530 199 1532 201
rect 1586 206 1588 208
rect 1580 196 1582 198
rect 1627 199 1629 201
rect 1675 199 1677 201
rect 1699 206 1701 208
rect 1705 196 1707 198
rect 1755 199 1757 201
rect 1765 199 1767 201
rect 1787 199 1789 201
rect 1797 199 1799 201
rect 1853 206 1855 208
rect 1847 196 1849 198
rect 1894 199 1896 201
rect 1985 206 1987 208
rect 1951 199 1953 201
rect 1961 198 1963 200
rect 1991 196 1993 198
rect 2041 199 2043 201
rect 2051 199 2053 201
rect 2073 199 2075 201
rect 2083 199 2085 201
rect 2139 206 2141 208
rect 2133 196 2135 198
rect 2180 199 2182 201
rect 2231 205 2233 207
rect 2249 204 2251 206
rect 2224 189 2226 191
rect 2299 205 2301 207
rect 2317 204 2319 206
rect 2292 189 2294 191
rect 33 119 35 121
rect 73 119 75 121
rect 103 122 105 124
rect 97 112 99 114
rect 153 119 155 121
rect 163 119 165 121
rect 185 119 187 121
rect 195 119 197 121
rect 245 122 247 124
rect 292 119 294 121
rect 251 112 253 114
rect 340 119 342 121
rect 370 122 372 124
rect 364 112 366 114
rect 420 119 422 121
rect 430 119 432 121
rect 452 119 454 121
rect 462 119 464 121
rect 512 122 514 124
rect 559 119 561 121
rect 518 112 520 114
rect 607 119 609 121
rect 637 122 639 124
rect 631 112 633 114
rect 687 119 689 121
rect 697 119 699 121
rect 719 119 721 121
rect 729 119 731 121
rect 779 122 781 124
rect 826 119 828 121
rect 785 112 787 114
rect 874 119 876 121
rect 904 122 906 124
rect 898 112 900 114
rect 954 119 956 121
rect 964 119 966 121
rect 986 119 988 121
rect 996 119 998 121
rect 1046 122 1048 124
rect 1093 119 1095 121
rect 1052 112 1054 114
rect 1141 119 1143 121
rect 1171 122 1173 124
rect 1165 112 1167 114
rect 1221 119 1223 121
rect 1231 119 1233 121
rect 1253 119 1255 121
rect 1263 119 1265 121
rect 1313 122 1315 124
rect 1360 119 1362 121
rect 1319 112 1321 114
rect 1408 119 1410 121
rect 1438 122 1440 124
rect 1432 112 1434 114
rect 1488 119 1490 121
rect 1498 119 1500 121
rect 1520 119 1522 121
rect 1530 119 1532 121
rect 1580 122 1582 124
rect 1627 119 1629 121
rect 1586 112 1588 114
rect 1675 119 1677 121
rect 1705 122 1707 124
rect 1699 112 1701 114
rect 1755 119 1757 121
rect 1765 119 1767 121
rect 1787 119 1789 121
rect 1797 119 1799 121
rect 1847 122 1849 124
rect 1894 119 1896 121
rect 1951 119 1953 121
rect 1961 120 1963 122
rect 1853 112 1855 114
rect 1991 122 1993 124
rect 1985 112 1987 114
rect 2041 119 2043 121
rect 2051 119 2053 121
rect 2073 119 2075 121
rect 2083 119 2085 121
rect 2133 122 2135 124
rect 2180 119 2182 121
rect 2139 112 2141 114
rect 2224 129 2226 131
rect 2231 113 2233 115
rect 2249 114 2251 116
rect 2292 129 2294 131
rect 2299 113 2301 115
rect 2317 114 2319 116
rect 33 55 35 57
rect 73 55 75 57
rect 97 62 99 64
rect 103 52 105 54
rect 153 55 155 57
rect 163 55 165 57
rect 185 55 187 57
rect 195 55 197 57
rect 251 62 253 64
rect 245 52 247 54
rect 292 55 294 57
rect 340 55 342 57
rect 364 62 366 64
rect 370 52 372 54
rect 420 55 422 57
rect 430 55 432 57
rect 452 55 454 57
rect 462 55 464 57
rect 518 62 520 64
rect 512 52 514 54
rect 559 55 561 57
rect 607 55 609 57
rect 631 62 633 64
rect 637 52 639 54
rect 687 55 689 57
rect 697 55 699 57
rect 719 55 721 57
rect 729 55 731 57
rect 785 62 787 64
rect 779 52 781 54
rect 826 55 828 57
rect 874 55 876 57
rect 898 62 900 64
rect 904 52 906 54
rect 954 55 956 57
rect 964 55 966 57
rect 986 55 988 57
rect 996 55 998 57
rect 1052 62 1054 64
rect 1046 52 1048 54
rect 1093 55 1095 57
rect 1141 55 1143 57
rect 1165 62 1167 64
rect 1171 52 1173 54
rect 1221 55 1223 57
rect 1231 55 1233 57
rect 1253 55 1255 57
rect 1263 55 1265 57
rect 1319 62 1321 64
rect 1313 52 1315 54
rect 1360 55 1362 57
rect 1408 55 1410 57
rect 1432 62 1434 64
rect 1438 52 1440 54
rect 1488 55 1490 57
rect 1498 55 1500 57
rect 1520 55 1522 57
rect 1530 55 1532 57
rect 1586 62 1588 64
rect 1580 52 1582 54
rect 1627 55 1629 57
rect 1675 55 1677 57
rect 1699 62 1701 64
rect 1705 52 1707 54
rect 1755 55 1757 57
rect 1765 55 1767 57
rect 1787 55 1789 57
rect 1797 55 1799 57
rect 1853 62 1855 64
rect 1847 52 1849 54
rect 1894 55 1896 57
rect 1985 62 1987 64
rect 1951 55 1953 57
rect 1961 54 1963 56
rect 1991 52 1993 54
rect 2041 55 2043 57
rect 2051 55 2053 57
rect 2073 55 2075 57
rect 2083 55 2085 57
rect 2139 62 2141 64
rect 2133 52 2135 54
rect 2180 55 2182 57
rect 2231 61 2233 63
rect 2249 60 2251 62
rect 2224 45 2226 47
rect 2299 61 2301 63
rect 2317 60 2319 62
rect 2292 45 2294 47
rect 33 -25 35 -23
rect 73 -25 75 -23
rect 103 -22 105 -20
rect 97 -32 99 -30
rect 153 -25 155 -23
rect 163 -25 165 -23
rect 185 -25 187 -23
rect 195 -25 197 -23
rect 245 -22 247 -20
rect 292 -25 294 -23
rect 251 -32 253 -30
rect 340 -25 342 -23
rect 370 -22 372 -20
rect 364 -32 366 -30
rect 420 -25 422 -23
rect 430 -25 432 -23
rect 452 -25 454 -23
rect 462 -25 464 -23
rect 512 -22 514 -20
rect 559 -25 561 -23
rect 518 -32 520 -30
rect 607 -25 609 -23
rect 637 -22 639 -20
rect 631 -32 633 -30
rect 687 -25 689 -23
rect 697 -25 699 -23
rect 719 -25 721 -23
rect 729 -25 731 -23
rect 779 -22 781 -20
rect 826 -25 828 -23
rect 785 -32 787 -30
rect 874 -25 876 -23
rect 904 -22 906 -20
rect 898 -32 900 -30
rect 954 -25 956 -23
rect 964 -25 966 -23
rect 986 -25 988 -23
rect 996 -25 998 -23
rect 1046 -22 1048 -20
rect 1093 -25 1095 -23
rect 1052 -32 1054 -30
rect 1141 -25 1143 -23
rect 1171 -22 1173 -20
rect 1165 -32 1167 -30
rect 1221 -25 1223 -23
rect 1231 -25 1233 -23
rect 1253 -25 1255 -23
rect 1263 -25 1265 -23
rect 1313 -22 1315 -20
rect 1360 -25 1362 -23
rect 1319 -32 1321 -30
rect 1408 -25 1410 -23
rect 1438 -22 1440 -20
rect 1432 -32 1434 -30
rect 1488 -25 1490 -23
rect 1498 -25 1500 -23
rect 1520 -25 1522 -23
rect 1530 -25 1532 -23
rect 1580 -22 1582 -20
rect 1627 -25 1629 -23
rect 1586 -32 1588 -30
rect 1675 -25 1677 -23
rect 1705 -22 1707 -20
rect 1699 -32 1701 -30
rect 1755 -25 1757 -23
rect 1765 -25 1767 -23
rect 1787 -25 1789 -23
rect 1797 -25 1799 -23
rect 1847 -22 1849 -20
rect 1894 -25 1896 -23
rect 1951 -25 1953 -23
rect 1961 -24 1963 -22
rect 1853 -32 1855 -30
rect 1991 -22 1993 -20
rect 1985 -32 1987 -30
rect 2041 -25 2043 -23
rect 2051 -25 2053 -23
rect 2073 -25 2075 -23
rect 2083 -25 2085 -23
rect 2133 -22 2135 -20
rect 2180 -25 2182 -23
rect 2139 -32 2141 -30
rect 2224 -15 2226 -13
rect 2231 -31 2233 -29
rect 2249 -30 2251 -28
rect 2292 -15 2294 -13
rect 2299 -31 2301 -29
rect 2317 -30 2319 -28
rect 33 -89 35 -87
rect 73 -89 75 -87
rect 97 -82 99 -80
rect 103 -92 105 -90
rect 153 -89 155 -87
rect 163 -89 165 -87
rect 185 -89 187 -87
rect 195 -89 197 -87
rect 251 -82 253 -80
rect 245 -92 247 -90
rect 292 -89 294 -87
rect 340 -89 342 -87
rect 364 -82 366 -80
rect 370 -92 372 -90
rect 420 -89 422 -87
rect 430 -89 432 -87
rect 452 -89 454 -87
rect 462 -89 464 -87
rect 518 -82 520 -80
rect 512 -92 514 -90
rect 559 -89 561 -87
rect 607 -89 609 -87
rect 631 -82 633 -80
rect 637 -92 639 -90
rect 687 -89 689 -87
rect 697 -89 699 -87
rect 719 -89 721 -87
rect 729 -89 731 -87
rect 785 -82 787 -80
rect 779 -92 781 -90
rect 826 -89 828 -87
rect 874 -89 876 -87
rect 898 -82 900 -80
rect 904 -92 906 -90
rect 954 -89 956 -87
rect 964 -89 966 -87
rect 986 -89 988 -87
rect 996 -89 998 -87
rect 1052 -82 1054 -80
rect 1046 -92 1048 -90
rect 1093 -89 1095 -87
rect 1141 -89 1143 -87
rect 1165 -82 1167 -80
rect 1171 -92 1173 -90
rect 1221 -89 1223 -87
rect 1231 -89 1233 -87
rect 1253 -89 1255 -87
rect 1263 -89 1265 -87
rect 1319 -82 1321 -80
rect 1313 -92 1315 -90
rect 1360 -89 1362 -87
rect 1408 -89 1410 -87
rect 1432 -82 1434 -80
rect 1438 -92 1440 -90
rect 1488 -89 1490 -87
rect 1498 -89 1500 -87
rect 1520 -89 1522 -87
rect 1530 -89 1532 -87
rect 1586 -82 1588 -80
rect 1580 -92 1582 -90
rect 1627 -89 1629 -87
rect 1675 -89 1677 -87
rect 1699 -82 1701 -80
rect 1705 -92 1707 -90
rect 1755 -89 1757 -87
rect 1765 -89 1767 -87
rect 1787 -89 1789 -87
rect 1797 -89 1799 -87
rect 1853 -82 1855 -80
rect 1847 -92 1849 -90
rect 1894 -89 1896 -87
rect 1985 -82 1987 -80
rect 1951 -89 1953 -87
rect 1961 -90 1963 -88
rect 1991 -92 1993 -90
rect 2041 -89 2043 -87
rect 2051 -89 2053 -87
rect 2073 -89 2075 -87
rect 2083 -89 2085 -87
rect 2139 -82 2141 -80
rect 2133 -92 2135 -90
rect 2180 -89 2182 -87
rect 2231 -83 2233 -81
rect 2249 -84 2251 -82
rect 2224 -99 2226 -97
rect 2299 -83 2301 -81
rect 2317 -84 2319 -82
rect 2292 -99 2294 -97
rect 33 -169 35 -167
rect 73 -169 75 -167
rect 103 -166 105 -164
rect 97 -176 99 -174
rect 153 -169 155 -167
rect 163 -169 165 -167
rect 185 -169 187 -167
rect 195 -169 197 -167
rect 245 -166 247 -164
rect 292 -169 294 -167
rect 251 -176 253 -174
rect 340 -169 342 -167
rect 370 -166 372 -164
rect 364 -176 366 -174
rect 420 -169 422 -167
rect 430 -169 432 -167
rect 452 -169 454 -167
rect 462 -169 464 -167
rect 512 -166 514 -164
rect 559 -169 561 -167
rect 518 -176 520 -174
rect 607 -169 609 -167
rect 637 -166 639 -164
rect 631 -176 633 -174
rect 687 -169 689 -167
rect 697 -169 699 -167
rect 719 -169 721 -167
rect 729 -169 731 -167
rect 779 -166 781 -164
rect 826 -169 828 -167
rect 785 -176 787 -174
rect 874 -169 876 -167
rect 904 -166 906 -164
rect 898 -176 900 -174
rect 954 -169 956 -167
rect 964 -169 966 -167
rect 986 -169 988 -167
rect 996 -169 998 -167
rect 1046 -166 1048 -164
rect 1093 -169 1095 -167
rect 1052 -176 1054 -174
rect 1141 -169 1143 -167
rect 1171 -166 1173 -164
rect 1165 -176 1167 -174
rect 1221 -169 1223 -167
rect 1231 -169 1233 -167
rect 1253 -169 1255 -167
rect 1263 -169 1265 -167
rect 1313 -166 1315 -164
rect 1360 -169 1362 -167
rect 1319 -176 1321 -174
rect 1408 -169 1410 -167
rect 1438 -166 1440 -164
rect 1432 -176 1434 -174
rect 1488 -169 1490 -167
rect 1498 -169 1500 -167
rect 1520 -169 1522 -167
rect 1530 -169 1532 -167
rect 1580 -166 1582 -164
rect 1627 -169 1629 -167
rect 1586 -176 1588 -174
rect 1675 -169 1677 -167
rect 1705 -166 1707 -164
rect 1699 -176 1701 -174
rect 1755 -169 1757 -167
rect 1765 -169 1767 -167
rect 1787 -169 1789 -167
rect 1797 -169 1799 -167
rect 1847 -166 1849 -164
rect 1894 -169 1896 -167
rect 1951 -169 1953 -167
rect 1961 -168 1963 -166
rect 1853 -176 1855 -174
rect 1991 -166 1993 -164
rect 1985 -176 1987 -174
rect 2041 -169 2043 -167
rect 2051 -169 2053 -167
rect 2073 -169 2075 -167
rect 2083 -169 2085 -167
rect 2133 -166 2135 -164
rect 2180 -169 2182 -167
rect 2139 -176 2141 -174
rect 2224 -159 2226 -157
rect 2231 -175 2233 -173
rect 2249 -174 2251 -172
rect 2292 -159 2294 -157
rect 2299 -175 2301 -173
rect 2317 -174 2319 -172
rect 33 -233 35 -231
rect 73 -233 75 -231
rect 97 -226 99 -224
rect 103 -236 105 -234
rect 153 -233 155 -231
rect 163 -233 165 -231
rect 185 -233 187 -231
rect 195 -233 197 -231
rect 251 -226 253 -224
rect 245 -236 247 -234
rect 292 -233 294 -231
rect 340 -233 342 -231
rect 364 -226 366 -224
rect 370 -236 372 -234
rect 420 -233 422 -231
rect 430 -233 432 -231
rect 452 -233 454 -231
rect 462 -233 464 -231
rect 518 -226 520 -224
rect 512 -236 514 -234
rect 559 -233 561 -231
rect 607 -233 609 -231
rect 631 -226 633 -224
rect 637 -236 639 -234
rect 687 -233 689 -231
rect 697 -233 699 -231
rect 719 -233 721 -231
rect 729 -233 731 -231
rect 785 -226 787 -224
rect 779 -236 781 -234
rect 826 -233 828 -231
rect 874 -233 876 -231
rect 898 -226 900 -224
rect 904 -236 906 -234
rect 954 -233 956 -231
rect 964 -233 966 -231
rect 986 -233 988 -231
rect 996 -233 998 -231
rect 1052 -226 1054 -224
rect 1046 -236 1048 -234
rect 1093 -233 1095 -231
rect 1141 -233 1143 -231
rect 1165 -226 1167 -224
rect 1171 -236 1173 -234
rect 1221 -233 1223 -231
rect 1231 -233 1233 -231
rect 1253 -233 1255 -231
rect 1263 -233 1265 -231
rect 1319 -226 1321 -224
rect 1313 -236 1315 -234
rect 1360 -233 1362 -231
rect 1408 -233 1410 -231
rect 1432 -226 1434 -224
rect 1438 -236 1440 -234
rect 1488 -233 1490 -231
rect 1498 -233 1500 -231
rect 1520 -233 1522 -231
rect 1530 -233 1532 -231
rect 1586 -226 1588 -224
rect 1580 -236 1582 -234
rect 1627 -233 1629 -231
rect 1675 -233 1677 -231
rect 1699 -226 1701 -224
rect 1705 -236 1707 -234
rect 1755 -233 1757 -231
rect 1765 -233 1767 -231
rect 1787 -233 1789 -231
rect 1797 -233 1799 -231
rect 1853 -226 1855 -224
rect 1847 -236 1849 -234
rect 1894 -233 1896 -231
rect 1985 -226 1987 -224
rect 1951 -233 1953 -231
rect 1961 -234 1963 -232
rect 1991 -236 1993 -234
rect 2041 -233 2043 -231
rect 2051 -233 2053 -231
rect 2073 -233 2075 -231
rect 2083 -233 2085 -231
rect 2139 -226 2141 -224
rect 2133 -236 2135 -234
rect 2180 -233 2182 -231
rect 2231 -227 2233 -225
rect 2249 -228 2251 -226
rect 2224 -243 2226 -241
rect 2299 -227 2301 -225
rect 2317 -228 2319 -226
rect 2292 -243 2294 -241
<< polyct1 >>
rect 13 271 15 273
rect 53 271 55 273
rect 23 263 25 265
rect 63 263 65 265
rect 117 263 119 265
rect 136 263 138 265
rect 143 263 145 265
rect 205 263 207 265
rect 212 263 214 265
rect 231 263 233 265
rect 272 270 274 272
rect 320 271 322 273
rect 282 263 284 265
rect 330 263 332 265
rect 384 263 386 265
rect 403 263 405 265
rect 410 263 412 265
rect 472 263 474 265
rect 479 263 481 265
rect 498 263 500 265
rect 539 270 541 272
rect 587 271 589 273
rect 549 263 551 265
rect 597 263 599 265
rect 651 263 653 265
rect 670 263 672 265
rect 677 263 679 265
rect 739 263 741 265
rect 746 263 748 265
rect 765 263 767 265
rect 806 270 808 272
rect 854 271 856 273
rect 816 263 818 265
rect 864 263 866 265
rect 918 263 920 265
rect 937 263 939 265
rect 944 263 946 265
rect 1006 263 1008 265
rect 1013 263 1015 265
rect 1032 263 1034 265
rect 1073 270 1075 272
rect 1121 271 1123 273
rect 1083 263 1085 265
rect 1131 263 1133 265
rect 1185 263 1187 265
rect 1204 263 1206 265
rect 1211 263 1213 265
rect 1273 263 1275 265
rect 1280 263 1282 265
rect 1299 263 1301 265
rect 1340 270 1342 272
rect 1388 271 1390 273
rect 1350 263 1352 265
rect 1398 263 1400 265
rect 1452 263 1454 265
rect 1471 263 1473 265
rect 1478 263 1480 265
rect 1540 263 1542 265
rect 1547 263 1549 265
rect 1566 263 1568 265
rect 1607 270 1609 272
rect 1655 271 1657 273
rect 1617 263 1619 265
rect 1665 263 1667 265
rect 1719 263 1721 265
rect 1738 263 1740 265
rect 1745 263 1747 265
rect 1807 263 1809 265
rect 1814 263 1816 265
rect 1833 263 1835 265
rect 1874 270 1876 272
rect 1914 271 1916 273
rect 1884 263 1886 265
rect 1930 258 1932 260
rect 2005 263 2007 265
rect 2024 263 2026 265
rect 2031 263 2033 265
rect 2093 263 2095 265
rect 2100 263 2102 265
rect 2119 263 2121 265
rect 2160 270 2162 272
rect 2201 283 2203 285
rect 2170 263 2172 265
rect 2269 283 2271 285
rect 2214 263 2216 265
rect 2241 268 2243 270
rect 2282 263 2284 265
rect 2309 268 2311 270
rect 23 199 25 201
rect 13 191 15 193
rect 63 199 65 201
rect 53 191 55 193
rect 117 199 119 201
rect 136 199 138 201
rect 143 199 145 201
rect 205 199 207 201
rect 212 199 214 201
rect 231 199 233 201
rect 282 199 284 201
rect 272 192 274 194
rect 330 199 332 201
rect 320 191 322 193
rect 384 199 386 201
rect 403 199 405 201
rect 410 199 412 201
rect 472 199 474 201
rect 479 199 481 201
rect 498 199 500 201
rect 549 199 551 201
rect 539 192 541 194
rect 597 199 599 201
rect 587 191 589 193
rect 651 199 653 201
rect 670 199 672 201
rect 677 199 679 201
rect 739 199 741 201
rect 746 199 748 201
rect 765 199 767 201
rect 816 199 818 201
rect 806 192 808 194
rect 864 199 866 201
rect 854 191 856 193
rect 918 199 920 201
rect 937 199 939 201
rect 944 199 946 201
rect 1006 199 1008 201
rect 1013 199 1015 201
rect 1032 199 1034 201
rect 1083 199 1085 201
rect 1073 192 1075 194
rect 1131 199 1133 201
rect 1121 191 1123 193
rect 1185 199 1187 201
rect 1204 199 1206 201
rect 1211 199 1213 201
rect 1273 199 1275 201
rect 1280 199 1282 201
rect 1299 199 1301 201
rect 1350 199 1352 201
rect 1340 192 1342 194
rect 1398 199 1400 201
rect 1388 191 1390 193
rect 1452 199 1454 201
rect 1471 199 1473 201
rect 1478 199 1480 201
rect 1540 199 1542 201
rect 1547 199 1549 201
rect 1566 199 1568 201
rect 1617 199 1619 201
rect 1607 192 1609 194
rect 1665 199 1667 201
rect 1655 191 1657 193
rect 1719 199 1721 201
rect 1738 199 1740 201
rect 1745 199 1747 201
rect 1807 199 1809 201
rect 1814 199 1816 201
rect 1833 199 1835 201
rect 1884 199 1886 201
rect 1930 204 1932 206
rect 1874 192 1876 194
rect 1914 191 1916 193
rect 2005 199 2007 201
rect 2024 199 2026 201
rect 2031 199 2033 201
rect 2093 199 2095 201
rect 2100 199 2102 201
rect 2119 199 2121 201
rect 2170 199 2172 201
rect 2160 192 2162 194
rect 2214 199 2216 201
rect 2241 194 2243 196
rect 2282 199 2284 201
rect 2201 179 2203 181
rect 2309 194 2311 196
rect 2269 179 2271 181
rect 13 127 15 129
rect 53 127 55 129
rect 23 119 25 121
rect 63 119 65 121
rect 117 119 119 121
rect 136 119 138 121
rect 143 119 145 121
rect 205 119 207 121
rect 212 119 214 121
rect 231 119 233 121
rect 272 126 274 128
rect 320 127 322 129
rect 282 119 284 121
rect 330 119 332 121
rect 384 119 386 121
rect 403 119 405 121
rect 410 119 412 121
rect 472 119 474 121
rect 479 119 481 121
rect 498 119 500 121
rect 539 126 541 128
rect 587 127 589 129
rect 549 119 551 121
rect 597 119 599 121
rect 651 119 653 121
rect 670 119 672 121
rect 677 119 679 121
rect 739 119 741 121
rect 746 119 748 121
rect 765 119 767 121
rect 806 126 808 128
rect 854 127 856 129
rect 816 119 818 121
rect 864 119 866 121
rect 918 119 920 121
rect 937 119 939 121
rect 944 119 946 121
rect 1006 119 1008 121
rect 1013 119 1015 121
rect 1032 119 1034 121
rect 1073 126 1075 128
rect 1121 127 1123 129
rect 1083 119 1085 121
rect 1131 119 1133 121
rect 1185 119 1187 121
rect 1204 119 1206 121
rect 1211 119 1213 121
rect 1273 119 1275 121
rect 1280 119 1282 121
rect 1299 119 1301 121
rect 1340 126 1342 128
rect 1388 127 1390 129
rect 1350 119 1352 121
rect 1398 119 1400 121
rect 1452 119 1454 121
rect 1471 119 1473 121
rect 1478 119 1480 121
rect 1540 119 1542 121
rect 1547 119 1549 121
rect 1566 119 1568 121
rect 1607 126 1609 128
rect 1655 127 1657 129
rect 1617 119 1619 121
rect 1665 119 1667 121
rect 1719 119 1721 121
rect 1738 119 1740 121
rect 1745 119 1747 121
rect 1807 119 1809 121
rect 1814 119 1816 121
rect 1833 119 1835 121
rect 1874 126 1876 128
rect 1914 127 1916 129
rect 1884 119 1886 121
rect 1930 114 1932 116
rect 2005 119 2007 121
rect 2024 119 2026 121
rect 2031 119 2033 121
rect 2093 119 2095 121
rect 2100 119 2102 121
rect 2119 119 2121 121
rect 2160 126 2162 128
rect 2201 139 2203 141
rect 2170 119 2172 121
rect 2269 139 2271 141
rect 2214 119 2216 121
rect 2241 124 2243 126
rect 2282 119 2284 121
rect 2309 124 2311 126
rect 23 55 25 57
rect 13 47 15 49
rect 63 55 65 57
rect 53 47 55 49
rect 117 55 119 57
rect 136 55 138 57
rect 143 55 145 57
rect 205 55 207 57
rect 212 55 214 57
rect 231 55 233 57
rect 282 55 284 57
rect 272 48 274 50
rect 330 55 332 57
rect 320 47 322 49
rect 384 55 386 57
rect 403 55 405 57
rect 410 55 412 57
rect 472 55 474 57
rect 479 55 481 57
rect 498 55 500 57
rect 549 55 551 57
rect 539 48 541 50
rect 597 55 599 57
rect 587 47 589 49
rect 651 55 653 57
rect 670 55 672 57
rect 677 55 679 57
rect 739 55 741 57
rect 746 55 748 57
rect 765 55 767 57
rect 816 55 818 57
rect 806 48 808 50
rect 864 55 866 57
rect 854 47 856 49
rect 918 55 920 57
rect 937 55 939 57
rect 944 55 946 57
rect 1006 55 1008 57
rect 1013 55 1015 57
rect 1032 55 1034 57
rect 1083 55 1085 57
rect 1073 48 1075 50
rect 1131 55 1133 57
rect 1121 47 1123 49
rect 1185 55 1187 57
rect 1204 55 1206 57
rect 1211 55 1213 57
rect 1273 55 1275 57
rect 1280 55 1282 57
rect 1299 55 1301 57
rect 1350 55 1352 57
rect 1340 48 1342 50
rect 1398 55 1400 57
rect 1388 47 1390 49
rect 1452 55 1454 57
rect 1471 55 1473 57
rect 1478 55 1480 57
rect 1540 55 1542 57
rect 1547 55 1549 57
rect 1566 55 1568 57
rect 1617 55 1619 57
rect 1607 48 1609 50
rect 1665 55 1667 57
rect 1655 47 1657 49
rect 1719 55 1721 57
rect 1738 55 1740 57
rect 1745 55 1747 57
rect 1807 55 1809 57
rect 1814 55 1816 57
rect 1833 55 1835 57
rect 1884 55 1886 57
rect 1930 60 1932 62
rect 1874 48 1876 50
rect 1914 47 1916 49
rect 2005 55 2007 57
rect 2024 55 2026 57
rect 2031 55 2033 57
rect 2093 55 2095 57
rect 2100 55 2102 57
rect 2119 55 2121 57
rect 2170 55 2172 57
rect 2160 48 2162 50
rect 2214 55 2216 57
rect 2241 50 2243 52
rect 2282 55 2284 57
rect 2201 35 2203 37
rect 2309 50 2311 52
rect 2269 35 2271 37
rect 13 -17 15 -15
rect 53 -17 55 -15
rect 23 -25 25 -23
rect 63 -25 65 -23
rect 117 -25 119 -23
rect 136 -25 138 -23
rect 143 -25 145 -23
rect 205 -25 207 -23
rect 212 -25 214 -23
rect 231 -25 233 -23
rect 272 -18 274 -16
rect 320 -17 322 -15
rect 282 -25 284 -23
rect 330 -25 332 -23
rect 384 -25 386 -23
rect 403 -25 405 -23
rect 410 -25 412 -23
rect 472 -25 474 -23
rect 479 -25 481 -23
rect 498 -25 500 -23
rect 539 -18 541 -16
rect 587 -17 589 -15
rect 549 -25 551 -23
rect 597 -25 599 -23
rect 651 -25 653 -23
rect 670 -25 672 -23
rect 677 -25 679 -23
rect 739 -25 741 -23
rect 746 -25 748 -23
rect 765 -25 767 -23
rect 806 -18 808 -16
rect 854 -17 856 -15
rect 816 -25 818 -23
rect 864 -25 866 -23
rect 918 -25 920 -23
rect 937 -25 939 -23
rect 944 -25 946 -23
rect 1006 -25 1008 -23
rect 1013 -25 1015 -23
rect 1032 -25 1034 -23
rect 1073 -18 1075 -16
rect 1121 -17 1123 -15
rect 1083 -25 1085 -23
rect 1131 -25 1133 -23
rect 1185 -25 1187 -23
rect 1204 -25 1206 -23
rect 1211 -25 1213 -23
rect 1273 -25 1275 -23
rect 1280 -25 1282 -23
rect 1299 -25 1301 -23
rect 1340 -18 1342 -16
rect 1388 -17 1390 -15
rect 1350 -25 1352 -23
rect 1398 -25 1400 -23
rect 1452 -25 1454 -23
rect 1471 -25 1473 -23
rect 1478 -25 1480 -23
rect 1540 -25 1542 -23
rect 1547 -25 1549 -23
rect 1566 -25 1568 -23
rect 1607 -18 1609 -16
rect 1655 -17 1657 -15
rect 1617 -25 1619 -23
rect 1665 -25 1667 -23
rect 1719 -25 1721 -23
rect 1738 -25 1740 -23
rect 1745 -25 1747 -23
rect 1807 -25 1809 -23
rect 1814 -25 1816 -23
rect 1833 -25 1835 -23
rect 1874 -18 1876 -16
rect 1914 -17 1916 -15
rect 1884 -25 1886 -23
rect 1930 -30 1932 -28
rect 2005 -25 2007 -23
rect 2024 -25 2026 -23
rect 2031 -25 2033 -23
rect 2093 -25 2095 -23
rect 2100 -25 2102 -23
rect 2119 -25 2121 -23
rect 2160 -18 2162 -16
rect 2201 -5 2203 -3
rect 2170 -25 2172 -23
rect 2269 -5 2271 -3
rect 2214 -25 2216 -23
rect 2241 -20 2243 -18
rect 2282 -25 2284 -23
rect 2309 -20 2311 -18
rect 23 -89 25 -87
rect 13 -97 15 -95
rect 63 -89 65 -87
rect 53 -97 55 -95
rect 117 -89 119 -87
rect 136 -89 138 -87
rect 143 -89 145 -87
rect 205 -89 207 -87
rect 212 -89 214 -87
rect 231 -89 233 -87
rect 282 -89 284 -87
rect 272 -96 274 -94
rect 330 -89 332 -87
rect 320 -97 322 -95
rect 384 -89 386 -87
rect 403 -89 405 -87
rect 410 -89 412 -87
rect 472 -89 474 -87
rect 479 -89 481 -87
rect 498 -89 500 -87
rect 549 -89 551 -87
rect 539 -96 541 -94
rect 597 -89 599 -87
rect 587 -97 589 -95
rect 651 -89 653 -87
rect 670 -89 672 -87
rect 677 -89 679 -87
rect 739 -89 741 -87
rect 746 -89 748 -87
rect 765 -89 767 -87
rect 816 -89 818 -87
rect 806 -96 808 -94
rect 864 -89 866 -87
rect 854 -97 856 -95
rect 918 -89 920 -87
rect 937 -89 939 -87
rect 944 -89 946 -87
rect 1006 -89 1008 -87
rect 1013 -89 1015 -87
rect 1032 -89 1034 -87
rect 1083 -89 1085 -87
rect 1073 -96 1075 -94
rect 1131 -89 1133 -87
rect 1121 -97 1123 -95
rect 1185 -89 1187 -87
rect 1204 -89 1206 -87
rect 1211 -89 1213 -87
rect 1273 -89 1275 -87
rect 1280 -89 1282 -87
rect 1299 -89 1301 -87
rect 1350 -89 1352 -87
rect 1340 -96 1342 -94
rect 1398 -89 1400 -87
rect 1388 -97 1390 -95
rect 1452 -89 1454 -87
rect 1471 -89 1473 -87
rect 1478 -89 1480 -87
rect 1540 -89 1542 -87
rect 1547 -89 1549 -87
rect 1566 -89 1568 -87
rect 1617 -89 1619 -87
rect 1607 -96 1609 -94
rect 1665 -89 1667 -87
rect 1655 -97 1657 -95
rect 1719 -89 1721 -87
rect 1738 -89 1740 -87
rect 1745 -89 1747 -87
rect 1807 -89 1809 -87
rect 1814 -89 1816 -87
rect 1833 -89 1835 -87
rect 1884 -89 1886 -87
rect 1930 -84 1932 -82
rect 1874 -96 1876 -94
rect 1914 -97 1916 -95
rect 2005 -89 2007 -87
rect 2024 -89 2026 -87
rect 2031 -89 2033 -87
rect 2093 -89 2095 -87
rect 2100 -89 2102 -87
rect 2119 -89 2121 -87
rect 2170 -89 2172 -87
rect 2160 -96 2162 -94
rect 2214 -89 2216 -87
rect 2241 -94 2243 -92
rect 2282 -89 2284 -87
rect 2201 -109 2203 -107
rect 2309 -94 2311 -92
rect 2269 -109 2271 -107
rect 13 -161 15 -159
rect 53 -161 55 -159
rect 23 -169 25 -167
rect 63 -169 65 -167
rect 117 -169 119 -167
rect 136 -169 138 -167
rect 143 -169 145 -167
rect 205 -169 207 -167
rect 212 -169 214 -167
rect 231 -169 233 -167
rect 272 -162 274 -160
rect 320 -161 322 -159
rect 282 -169 284 -167
rect 330 -169 332 -167
rect 384 -169 386 -167
rect 403 -169 405 -167
rect 410 -169 412 -167
rect 472 -169 474 -167
rect 479 -169 481 -167
rect 498 -169 500 -167
rect 539 -162 541 -160
rect 587 -161 589 -159
rect 549 -169 551 -167
rect 597 -169 599 -167
rect 651 -169 653 -167
rect 670 -169 672 -167
rect 677 -169 679 -167
rect 739 -169 741 -167
rect 746 -169 748 -167
rect 765 -169 767 -167
rect 806 -162 808 -160
rect 854 -161 856 -159
rect 816 -169 818 -167
rect 864 -169 866 -167
rect 918 -169 920 -167
rect 937 -169 939 -167
rect 944 -169 946 -167
rect 1006 -169 1008 -167
rect 1013 -169 1015 -167
rect 1032 -169 1034 -167
rect 1073 -162 1075 -160
rect 1121 -161 1123 -159
rect 1083 -169 1085 -167
rect 1131 -169 1133 -167
rect 1185 -169 1187 -167
rect 1204 -169 1206 -167
rect 1211 -169 1213 -167
rect 1273 -169 1275 -167
rect 1280 -169 1282 -167
rect 1299 -169 1301 -167
rect 1340 -162 1342 -160
rect 1388 -161 1390 -159
rect 1350 -169 1352 -167
rect 1398 -169 1400 -167
rect 1452 -169 1454 -167
rect 1471 -169 1473 -167
rect 1478 -169 1480 -167
rect 1540 -169 1542 -167
rect 1547 -169 1549 -167
rect 1566 -169 1568 -167
rect 1607 -162 1609 -160
rect 1655 -161 1657 -159
rect 1617 -169 1619 -167
rect 1665 -169 1667 -167
rect 1719 -169 1721 -167
rect 1738 -169 1740 -167
rect 1745 -169 1747 -167
rect 1807 -169 1809 -167
rect 1814 -169 1816 -167
rect 1833 -169 1835 -167
rect 1874 -162 1876 -160
rect 1914 -161 1916 -159
rect 1884 -169 1886 -167
rect 1930 -174 1932 -172
rect 2005 -169 2007 -167
rect 2024 -169 2026 -167
rect 2031 -169 2033 -167
rect 2093 -169 2095 -167
rect 2100 -169 2102 -167
rect 2119 -169 2121 -167
rect 2160 -162 2162 -160
rect 2201 -149 2203 -147
rect 2170 -169 2172 -167
rect 2269 -149 2271 -147
rect 2214 -169 2216 -167
rect 2241 -164 2243 -162
rect 2282 -169 2284 -167
rect 2309 -164 2311 -162
rect 23 -233 25 -231
rect 13 -241 15 -239
rect 63 -233 65 -231
rect 53 -241 55 -239
rect 117 -233 119 -231
rect 136 -233 138 -231
rect 143 -233 145 -231
rect 205 -233 207 -231
rect 212 -233 214 -231
rect 231 -233 233 -231
rect 282 -233 284 -231
rect 272 -240 274 -238
rect 330 -233 332 -231
rect 320 -241 322 -239
rect 384 -233 386 -231
rect 403 -233 405 -231
rect 410 -233 412 -231
rect 472 -233 474 -231
rect 479 -233 481 -231
rect 498 -233 500 -231
rect 549 -233 551 -231
rect 539 -240 541 -238
rect 597 -233 599 -231
rect 587 -241 589 -239
rect 651 -233 653 -231
rect 670 -233 672 -231
rect 677 -233 679 -231
rect 739 -233 741 -231
rect 746 -233 748 -231
rect 765 -233 767 -231
rect 816 -233 818 -231
rect 806 -240 808 -238
rect 864 -233 866 -231
rect 854 -241 856 -239
rect 918 -233 920 -231
rect 937 -233 939 -231
rect 944 -233 946 -231
rect 1006 -233 1008 -231
rect 1013 -233 1015 -231
rect 1032 -233 1034 -231
rect 1083 -233 1085 -231
rect 1073 -240 1075 -238
rect 1131 -233 1133 -231
rect 1121 -241 1123 -239
rect 1185 -233 1187 -231
rect 1204 -233 1206 -231
rect 1211 -233 1213 -231
rect 1273 -233 1275 -231
rect 1280 -233 1282 -231
rect 1299 -233 1301 -231
rect 1350 -233 1352 -231
rect 1340 -240 1342 -238
rect 1398 -233 1400 -231
rect 1388 -241 1390 -239
rect 1452 -233 1454 -231
rect 1471 -233 1473 -231
rect 1478 -233 1480 -231
rect 1540 -233 1542 -231
rect 1547 -233 1549 -231
rect 1566 -233 1568 -231
rect 1617 -233 1619 -231
rect 1607 -240 1609 -238
rect 1665 -233 1667 -231
rect 1655 -241 1657 -239
rect 1719 -233 1721 -231
rect 1738 -233 1740 -231
rect 1745 -233 1747 -231
rect 1807 -233 1809 -231
rect 1814 -233 1816 -231
rect 1833 -233 1835 -231
rect 1884 -233 1886 -231
rect 1930 -228 1932 -226
rect 1874 -240 1876 -238
rect 1914 -241 1916 -239
rect 2005 -233 2007 -231
rect 2024 -233 2026 -231
rect 2031 -233 2033 -231
rect 2093 -233 2095 -231
rect 2100 -233 2102 -231
rect 2119 -233 2121 -231
rect 2170 -233 2172 -231
rect 2160 -240 2162 -238
rect 2214 -233 2216 -231
rect 2241 -238 2243 -236
rect 2282 -233 2284 -231
rect 2201 -253 2203 -251
rect 2309 -238 2311 -236
rect 2269 -253 2271 -251
<< ndifct0 >>
rect 10 247 12 249
rect 50 247 52 249
rect 100 243 102 245
rect 110 246 112 248
rect 120 254 122 256
rect 130 254 132 256
rect 130 247 132 249
rect 140 247 142 249
rect 157 240 159 242
rect 191 240 193 242
rect 218 254 220 256
rect 208 247 210 249
rect 218 247 220 249
rect 228 254 230 256
rect 279 254 281 256
rect 238 246 240 248
rect 248 243 250 245
rect 269 241 271 243
rect 317 247 319 249
rect 288 241 290 243
rect 367 243 369 245
rect 377 246 379 248
rect 387 254 389 256
rect 397 254 399 256
rect 397 247 399 249
rect 407 247 409 249
rect 424 240 426 242
rect 458 240 460 242
rect 485 254 487 256
rect 475 247 477 249
rect 485 247 487 249
rect 495 254 497 256
rect 546 254 548 256
rect 505 246 507 248
rect 515 243 517 245
rect 536 241 538 243
rect 584 247 586 249
rect 555 241 557 243
rect 634 243 636 245
rect 644 246 646 248
rect 654 254 656 256
rect 664 254 666 256
rect 664 247 666 249
rect 674 247 676 249
rect 691 240 693 242
rect 725 240 727 242
rect 752 254 754 256
rect 742 247 744 249
rect 752 247 754 249
rect 762 254 764 256
rect 813 254 815 256
rect 772 246 774 248
rect 782 243 784 245
rect 803 241 805 243
rect 851 247 853 249
rect 822 241 824 243
rect 901 243 903 245
rect 911 246 913 248
rect 921 254 923 256
rect 931 254 933 256
rect 931 247 933 249
rect 941 247 943 249
rect 958 240 960 242
rect 992 240 994 242
rect 1019 254 1021 256
rect 1009 247 1011 249
rect 1019 247 1021 249
rect 1029 254 1031 256
rect 1080 254 1082 256
rect 1039 246 1041 248
rect 1049 243 1051 245
rect 1070 241 1072 243
rect 1118 247 1120 249
rect 1089 241 1091 243
rect 1168 243 1170 245
rect 1178 246 1180 248
rect 1188 254 1190 256
rect 1198 254 1200 256
rect 1198 247 1200 249
rect 1208 247 1210 249
rect 1225 240 1227 242
rect 1259 240 1261 242
rect 1286 254 1288 256
rect 1276 247 1278 249
rect 1286 247 1288 249
rect 1296 254 1298 256
rect 1347 254 1349 256
rect 1306 246 1308 248
rect 1316 243 1318 245
rect 1337 241 1339 243
rect 1385 247 1387 249
rect 1356 241 1358 243
rect 1435 243 1437 245
rect 1445 246 1447 248
rect 1455 254 1457 256
rect 1465 254 1467 256
rect 1465 247 1467 249
rect 1475 247 1477 249
rect 1492 240 1494 242
rect 1526 240 1528 242
rect 1553 254 1555 256
rect 1543 247 1545 249
rect 1553 247 1555 249
rect 1563 254 1565 256
rect 1614 254 1616 256
rect 1573 246 1575 248
rect 1583 243 1585 245
rect 1604 241 1606 243
rect 1652 247 1654 249
rect 1623 241 1625 243
rect 1702 243 1704 245
rect 1712 246 1714 248
rect 1722 254 1724 256
rect 1732 254 1734 256
rect 1732 247 1734 249
rect 1742 247 1744 249
rect 1759 240 1761 242
rect 1793 240 1795 242
rect 1820 254 1822 256
rect 1810 247 1812 249
rect 1820 247 1822 249
rect 1830 254 1832 256
rect 1881 254 1883 256
rect 1840 246 1842 248
rect 1850 243 1852 245
rect 1914 254 1916 256
rect 1871 241 1873 243
rect 1928 246 1930 248
rect 1940 249 1942 251
rect 1890 241 1892 243
rect 1988 243 1990 245
rect 1998 246 2000 248
rect 2008 254 2010 256
rect 2018 254 2020 256
rect 2018 247 2020 249
rect 2028 247 2030 249
rect 2045 240 2047 242
rect 2079 240 2081 242
rect 2106 254 2108 256
rect 2096 247 2098 249
rect 2106 247 2108 249
rect 2116 254 2118 256
rect 2167 254 2169 256
rect 2126 246 2128 248
rect 2136 243 2138 245
rect 2157 241 2159 243
rect 2201 248 2203 250
rect 2211 248 2213 250
rect 2176 241 2178 243
rect 2228 246 2230 248
rect 2245 246 2247 248
rect 2269 248 2271 250
rect 2279 248 2281 250
rect 2296 246 2298 248
rect 2313 246 2315 248
rect 10 215 12 217
rect 50 215 52 217
rect 100 219 102 221
rect 110 216 112 218
rect 120 208 122 210
rect 130 215 132 217
rect 140 215 142 217
rect 130 208 132 210
rect 157 222 159 224
rect 191 222 193 224
rect 208 215 210 217
rect 218 215 220 217
rect 218 208 220 210
rect 228 208 230 210
rect 238 216 240 218
rect 248 219 250 221
rect 269 221 271 223
rect 288 221 290 223
rect 317 215 319 217
rect 279 208 281 210
rect 367 219 369 221
rect 377 216 379 218
rect 387 208 389 210
rect 397 215 399 217
rect 407 215 409 217
rect 397 208 399 210
rect 424 222 426 224
rect 458 222 460 224
rect 475 215 477 217
rect 485 215 487 217
rect 485 208 487 210
rect 495 208 497 210
rect 505 216 507 218
rect 515 219 517 221
rect 536 221 538 223
rect 555 221 557 223
rect 584 215 586 217
rect 546 208 548 210
rect 634 219 636 221
rect 644 216 646 218
rect 654 208 656 210
rect 664 215 666 217
rect 674 215 676 217
rect 664 208 666 210
rect 691 222 693 224
rect 725 222 727 224
rect 742 215 744 217
rect 752 215 754 217
rect 752 208 754 210
rect 762 208 764 210
rect 772 216 774 218
rect 782 219 784 221
rect 803 221 805 223
rect 822 221 824 223
rect 851 215 853 217
rect 813 208 815 210
rect 901 219 903 221
rect 911 216 913 218
rect 921 208 923 210
rect 931 215 933 217
rect 941 215 943 217
rect 931 208 933 210
rect 958 222 960 224
rect 992 222 994 224
rect 1009 215 1011 217
rect 1019 215 1021 217
rect 1019 208 1021 210
rect 1029 208 1031 210
rect 1039 216 1041 218
rect 1049 219 1051 221
rect 1070 221 1072 223
rect 1089 221 1091 223
rect 1118 215 1120 217
rect 1080 208 1082 210
rect 1168 219 1170 221
rect 1178 216 1180 218
rect 1188 208 1190 210
rect 1198 215 1200 217
rect 1208 215 1210 217
rect 1198 208 1200 210
rect 1225 222 1227 224
rect 1259 222 1261 224
rect 1276 215 1278 217
rect 1286 215 1288 217
rect 1286 208 1288 210
rect 1296 208 1298 210
rect 1306 216 1308 218
rect 1316 219 1318 221
rect 1337 221 1339 223
rect 1356 221 1358 223
rect 1385 215 1387 217
rect 1347 208 1349 210
rect 1435 219 1437 221
rect 1445 216 1447 218
rect 1455 208 1457 210
rect 1465 215 1467 217
rect 1475 215 1477 217
rect 1465 208 1467 210
rect 1492 222 1494 224
rect 1526 222 1528 224
rect 1543 215 1545 217
rect 1553 215 1555 217
rect 1553 208 1555 210
rect 1563 208 1565 210
rect 1573 216 1575 218
rect 1583 219 1585 221
rect 1604 221 1606 223
rect 1623 221 1625 223
rect 1652 215 1654 217
rect 1614 208 1616 210
rect 1702 219 1704 221
rect 1712 216 1714 218
rect 1722 208 1724 210
rect 1732 215 1734 217
rect 1742 215 1744 217
rect 1732 208 1734 210
rect 1759 222 1761 224
rect 1793 222 1795 224
rect 1810 215 1812 217
rect 1820 215 1822 217
rect 1820 208 1822 210
rect 1830 208 1832 210
rect 1840 216 1842 218
rect 1850 219 1852 221
rect 1871 221 1873 223
rect 1890 221 1892 223
rect 1928 216 1930 218
rect 1881 208 1883 210
rect 1914 208 1916 210
rect 1940 213 1942 215
rect 1988 219 1990 221
rect 1998 216 2000 218
rect 2008 208 2010 210
rect 2018 215 2020 217
rect 2028 215 2030 217
rect 2018 208 2020 210
rect 2045 222 2047 224
rect 2079 222 2081 224
rect 2096 215 2098 217
rect 2106 215 2108 217
rect 2106 208 2108 210
rect 2116 208 2118 210
rect 2126 216 2128 218
rect 2136 219 2138 221
rect 2157 221 2159 223
rect 2176 221 2178 223
rect 2167 208 2169 210
rect 2201 214 2203 216
rect 2211 214 2213 216
rect 2228 216 2230 218
rect 2245 216 2247 218
rect 2269 214 2271 216
rect 2279 214 2281 216
rect 2296 216 2298 218
rect 2313 216 2315 218
rect 10 103 12 105
rect 50 103 52 105
rect 100 99 102 101
rect 110 102 112 104
rect 120 110 122 112
rect 130 110 132 112
rect 130 103 132 105
rect 140 103 142 105
rect 157 96 159 98
rect 191 96 193 98
rect 218 110 220 112
rect 208 103 210 105
rect 218 103 220 105
rect 228 110 230 112
rect 279 110 281 112
rect 238 102 240 104
rect 248 99 250 101
rect 269 97 271 99
rect 317 103 319 105
rect 288 97 290 99
rect 367 99 369 101
rect 377 102 379 104
rect 387 110 389 112
rect 397 110 399 112
rect 397 103 399 105
rect 407 103 409 105
rect 424 96 426 98
rect 458 96 460 98
rect 485 110 487 112
rect 475 103 477 105
rect 485 103 487 105
rect 495 110 497 112
rect 546 110 548 112
rect 505 102 507 104
rect 515 99 517 101
rect 536 97 538 99
rect 584 103 586 105
rect 555 97 557 99
rect 634 99 636 101
rect 644 102 646 104
rect 654 110 656 112
rect 664 110 666 112
rect 664 103 666 105
rect 674 103 676 105
rect 691 96 693 98
rect 725 96 727 98
rect 752 110 754 112
rect 742 103 744 105
rect 752 103 754 105
rect 762 110 764 112
rect 813 110 815 112
rect 772 102 774 104
rect 782 99 784 101
rect 803 97 805 99
rect 851 103 853 105
rect 822 97 824 99
rect 901 99 903 101
rect 911 102 913 104
rect 921 110 923 112
rect 931 110 933 112
rect 931 103 933 105
rect 941 103 943 105
rect 958 96 960 98
rect 992 96 994 98
rect 1019 110 1021 112
rect 1009 103 1011 105
rect 1019 103 1021 105
rect 1029 110 1031 112
rect 1080 110 1082 112
rect 1039 102 1041 104
rect 1049 99 1051 101
rect 1070 97 1072 99
rect 1118 103 1120 105
rect 1089 97 1091 99
rect 1168 99 1170 101
rect 1178 102 1180 104
rect 1188 110 1190 112
rect 1198 110 1200 112
rect 1198 103 1200 105
rect 1208 103 1210 105
rect 1225 96 1227 98
rect 1259 96 1261 98
rect 1286 110 1288 112
rect 1276 103 1278 105
rect 1286 103 1288 105
rect 1296 110 1298 112
rect 1347 110 1349 112
rect 1306 102 1308 104
rect 1316 99 1318 101
rect 1337 97 1339 99
rect 1385 103 1387 105
rect 1356 97 1358 99
rect 1435 99 1437 101
rect 1445 102 1447 104
rect 1455 110 1457 112
rect 1465 110 1467 112
rect 1465 103 1467 105
rect 1475 103 1477 105
rect 1492 96 1494 98
rect 1526 96 1528 98
rect 1553 110 1555 112
rect 1543 103 1545 105
rect 1553 103 1555 105
rect 1563 110 1565 112
rect 1614 110 1616 112
rect 1573 102 1575 104
rect 1583 99 1585 101
rect 1604 97 1606 99
rect 1652 103 1654 105
rect 1623 97 1625 99
rect 1702 99 1704 101
rect 1712 102 1714 104
rect 1722 110 1724 112
rect 1732 110 1734 112
rect 1732 103 1734 105
rect 1742 103 1744 105
rect 1759 96 1761 98
rect 1793 96 1795 98
rect 1820 110 1822 112
rect 1810 103 1812 105
rect 1820 103 1822 105
rect 1830 110 1832 112
rect 1881 110 1883 112
rect 1840 102 1842 104
rect 1850 99 1852 101
rect 1914 110 1916 112
rect 1871 97 1873 99
rect 1928 102 1930 104
rect 1940 105 1942 107
rect 1890 97 1892 99
rect 1988 99 1990 101
rect 1998 102 2000 104
rect 2008 110 2010 112
rect 2018 110 2020 112
rect 2018 103 2020 105
rect 2028 103 2030 105
rect 2045 96 2047 98
rect 2079 96 2081 98
rect 2106 110 2108 112
rect 2096 103 2098 105
rect 2106 103 2108 105
rect 2116 110 2118 112
rect 2167 110 2169 112
rect 2126 102 2128 104
rect 2136 99 2138 101
rect 2157 97 2159 99
rect 2201 104 2203 106
rect 2211 104 2213 106
rect 2176 97 2178 99
rect 2228 102 2230 104
rect 2245 102 2247 104
rect 2269 104 2271 106
rect 2279 104 2281 106
rect 2296 102 2298 104
rect 2313 102 2315 104
rect 10 71 12 73
rect 50 71 52 73
rect 100 75 102 77
rect 110 72 112 74
rect 120 64 122 66
rect 130 71 132 73
rect 140 71 142 73
rect 130 64 132 66
rect 157 78 159 80
rect 191 78 193 80
rect 208 71 210 73
rect 218 71 220 73
rect 218 64 220 66
rect 228 64 230 66
rect 238 72 240 74
rect 248 75 250 77
rect 269 77 271 79
rect 288 77 290 79
rect 317 71 319 73
rect 279 64 281 66
rect 367 75 369 77
rect 377 72 379 74
rect 387 64 389 66
rect 397 71 399 73
rect 407 71 409 73
rect 397 64 399 66
rect 424 78 426 80
rect 458 78 460 80
rect 475 71 477 73
rect 485 71 487 73
rect 485 64 487 66
rect 495 64 497 66
rect 505 72 507 74
rect 515 75 517 77
rect 536 77 538 79
rect 555 77 557 79
rect 584 71 586 73
rect 546 64 548 66
rect 634 75 636 77
rect 644 72 646 74
rect 654 64 656 66
rect 664 71 666 73
rect 674 71 676 73
rect 664 64 666 66
rect 691 78 693 80
rect 725 78 727 80
rect 742 71 744 73
rect 752 71 754 73
rect 752 64 754 66
rect 762 64 764 66
rect 772 72 774 74
rect 782 75 784 77
rect 803 77 805 79
rect 822 77 824 79
rect 851 71 853 73
rect 813 64 815 66
rect 901 75 903 77
rect 911 72 913 74
rect 921 64 923 66
rect 931 71 933 73
rect 941 71 943 73
rect 931 64 933 66
rect 958 78 960 80
rect 992 78 994 80
rect 1009 71 1011 73
rect 1019 71 1021 73
rect 1019 64 1021 66
rect 1029 64 1031 66
rect 1039 72 1041 74
rect 1049 75 1051 77
rect 1070 77 1072 79
rect 1089 77 1091 79
rect 1118 71 1120 73
rect 1080 64 1082 66
rect 1168 75 1170 77
rect 1178 72 1180 74
rect 1188 64 1190 66
rect 1198 71 1200 73
rect 1208 71 1210 73
rect 1198 64 1200 66
rect 1225 78 1227 80
rect 1259 78 1261 80
rect 1276 71 1278 73
rect 1286 71 1288 73
rect 1286 64 1288 66
rect 1296 64 1298 66
rect 1306 72 1308 74
rect 1316 75 1318 77
rect 1337 77 1339 79
rect 1356 77 1358 79
rect 1385 71 1387 73
rect 1347 64 1349 66
rect 1435 75 1437 77
rect 1445 72 1447 74
rect 1455 64 1457 66
rect 1465 71 1467 73
rect 1475 71 1477 73
rect 1465 64 1467 66
rect 1492 78 1494 80
rect 1526 78 1528 80
rect 1543 71 1545 73
rect 1553 71 1555 73
rect 1553 64 1555 66
rect 1563 64 1565 66
rect 1573 72 1575 74
rect 1583 75 1585 77
rect 1604 77 1606 79
rect 1623 77 1625 79
rect 1652 71 1654 73
rect 1614 64 1616 66
rect 1702 75 1704 77
rect 1712 72 1714 74
rect 1722 64 1724 66
rect 1732 71 1734 73
rect 1742 71 1744 73
rect 1732 64 1734 66
rect 1759 78 1761 80
rect 1793 78 1795 80
rect 1810 71 1812 73
rect 1820 71 1822 73
rect 1820 64 1822 66
rect 1830 64 1832 66
rect 1840 72 1842 74
rect 1850 75 1852 77
rect 1871 77 1873 79
rect 1890 77 1892 79
rect 1928 72 1930 74
rect 1881 64 1883 66
rect 1914 64 1916 66
rect 1940 69 1942 71
rect 1988 75 1990 77
rect 1998 72 2000 74
rect 2008 64 2010 66
rect 2018 71 2020 73
rect 2028 71 2030 73
rect 2018 64 2020 66
rect 2045 78 2047 80
rect 2079 78 2081 80
rect 2096 71 2098 73
rect 2106 71 2108 73
rect 2106 64 2108 66
rect 2116 64 2118 66
rect 2126 72 2128 74
rect 2136 75 2138 77
rect 2157 77 2159 79
rect 2176 77 2178 79
rect 2167 64 2169 66
rect 2201 70 2203 72
rect 2211 70 2213 72
rect 2228 72 2230 74
rect 2245 72 2247 74
rect 2269 70 2271 72
rect 2279 70 2281 72
rect 2296 72 2298 74
rect 2313 72 2315 74
rect 10 -41 12 -39
rect 50 -41 52 -39
rect 100 -45 102 -43
rect 110 -42 112 -40
rect 120 -34 122 -32
rect 130 -34 132 -32
rect 130 -41 132 -39
rect 140 -41 142 -39
rect 157 -48 159 -46
rect 191 -48 193 -46
rect 218 -34 220 -32
rect 208 -41 210 -39
rect 218 -41 220 -39
rect 228 -34 230 -32
rect 279 -34 281 -32
rect 238 -42 240 -40
rect 248 -45 250 -43
rect 269 -47 271 -45
rect 317 -41 319 -39
rect 288 -47 290 -45
rect 367 -45 369 -43
rect 377 -42 379 -40
rect 387 -34 389 -32
rect 397 -34 399 -32
rect 397 -41 399 -39
rect 407 -41 409 -39
rect 424 -48 426 -46
rect 458 -48 460 -46
rect 485 -34 487 -32
rect 475 -41 477 -39
rect 485 -41 487 -39
rect 495 -34 497 -32
rect 546 -34 548 -32
rect 505 -42 507 -40
rect 515 -45 517 -43
rect 536 -47 538 -45
rect 584 -41 586 -39
rect 555 -47 557 -45
rect 634 -45 636 -43
rect 644 -42 646 -40
rect 654 -34 656 -32
rect 664 -34 666 -32
rect 664 -41 666 -39
rect 674 -41 676 -39
rect 691 -48 693 -46
rect 725 -48 727 -46
rect 752 -34 754 -32
rect 742 -41 744 -39
rect 752 -41 754 -39
rect 762 -34 764 -32
rect 813 -34 815 -32
rect 772 -42 774 -40
rect 782 -45 784 -43
rect 803 -47 805 -45
rect 851 -41 853 -39
rect 822 -47 824 -45
rect 901 -45 903 -43
rect 911 -42 913 -40
rect 921 -34 923 -32
rect 931 -34 933 -32
rect 931 -41 933 -39
rect 941 -41 943 -39
rect 958 -48 960 -46
rect 992 -48 994 -46
rect 1019 -34 1021 -32
rect 1009 -41 1011 -39
rect 1019 -41 1021 -39
rect 1029 -34 1031 -32
rect 1080 -34 1082 -32
rect 1039 -42 1041 -40
rect 1049 -45 1051 -43
rect 1070 -47 1072 -45
rect 1118 -41 1120 -39
rect 1089 -47 1091 -45
rect 1168 -45 1170 -43
rect 1178 -42 1180 -40
rect 1188 -34 1190 -32
rect 1198 -34 1200 -32
rect 1198 -41 1200 -39
rect 1208 -41 1210 -39
rect 1225 -48 1227 -46
rect 1259 -48 1261 -46
rect 1286 -34 1288 -32
rect 1276 -41 1278 -39
rect 1286 -41 1288 -39
rect 1296 -34 1298 -32
rect 1347 -34 1349 -32
rect 1306 -42 1308 -40
rect 1316 -45 1318 -43
rect 1337 -47 1339 -45
rect 1385 -41 1387 -39
rect 1356 -47 1358 -45
rect 1435 -45 1437 -43
rect 1445 -42 1447 -40
rect 1455 -34 1457 -32
rect 1465 -34 1467 -32
rect 1465 -41 1467 -39
rect 1475 -41 1477 -39
rect 1492 -48 1494 -46
rect 1526 -48 1528 -46
rect 1553 -34 1555 -32
rect 1543 -41 1545 -39
rect 1553 -41 1555 -39
rect 1563 -34 1565 -32
rect 1614 -34 1616 -32
rect 1573 -42 1575 -40
rect 1583 -45 1585 -43
rect 1604 -47 1606 -45
rect 1652 -41 1654 -39
rect 1623 -47 1625 -45
rect 1702 -45 1704 -43
rect 1712 -42 1714 -40
rect 1722 -34 1724 -32
rect 1732 -34 1734 -32
rect 1732 -41 1734 -39
rect 1742 -41 1744 -39
rect 1759 -48 1761 -46
rect 1793 -48 1795 -46
rect 1820 -34 1822 -32
rect 1810 -41 1812 -39
rect 1820 -41 1822 -39
rect 1830 -34 1832 -32
rect 1881 -34 1883 -32
rect 1840 -42 1842 -40
rect 1850 -45 1852 -43
rect 1914 -34 1916 -32
rect 1871 -47 1873 -45
rect 1928 -42 1930 -40
rect 1940 -39 1942 -37
rect 1890 -47 1892 -45
rect 1988 -45 1990 -43
rect 1998 -42 2000 -40
rect 2008 -34 2010 -32
rect 2018 -34 2020 -32
rect 2018 -41 2020 -39
rect 2028 -41 2030 -39
rect 2045 -48 2047 -46
rect 2079 -48 2081 -46
rect 2106 -34 2108 -32
rect 2096 -41 2098 -39
rect 2106 -41 2108 -39
rect 2116 -34 2118 -32
rect 2167 -34 2169 -32
rect 2126 -42 2128 -40
rect 2136 -45 2138 -43
rect 2157 -47 2159 -45
rect 2201 -40 2203 -38
rect 2211 -40 2213 -38
rect 2176 -47 2178 -45
rect 2228 -42 2230 -40
rect 2245 -42 2247 -40
rect 2269 -40 2271 -38
rect 2279 -40 2281 -38
rect 2296 -42 2298 -40
rect 2313 -42 2315 -40
rect 10 -73 12 -71
rect 50 -73 52 -71
rect 100 -69 102 -67
rect 110 -72 112 -70
rect 120 -80 122 -78
rect 130 -73 132 -71
rect 140 -73 142 -71
rect 130 -80 132 -78
rect 157 -66 159 -64
rect 191 -66 193 -64
rect 208 -73 210 -71
rect 218 -73 220 -71
rect 218 -80 220 -78
rect 228 -80 230 -78
rect 238 -72 240 -70
rect 248 -69 250 -67
rect 269 -67 271 -65
rect 288 -67 290 -65
rect 317 -73 319 -71
rect 279 -80 281 -78
rect 367 -69 369 -67
rect 377 -72 379 -70
rect 387 -80 389 -78
rect 397 -73 399 -71
rect 407 -73 409 -71
rect 397 -80 399 -78
rect 424 -66 426 -64
rect 458 -66 460 -64
rect 475 -73 477 -71
rect 485 -73 487 -71
rect 485 -80 487 -78
rect 495 -80 497 -78
rect 505 -72 507 -70
rect 515 -69 517 -67
rect 536 -67 538 -65
rect 555 -67 557 -65
rect 584 -73 586 -71
rect 546 -80 548 -78
rect 634 -69 636 -67
rect 644 -72 646 -70
rect 654 -80 656 -78
rect 664 -73 666 -71
rect 674 -73 676 -71
rect 664 -80 666 -78
rect 691 -66 693 -64
rect 725 -66 727 -64
rect 742 -73 744 -71
rect 752 -73 754 -71
rect 752 -80 754 -78
rect 762 -80 764 -78
rect 772 -72 774 -70
rect 782 -69 784 -67
rect 803 -67 805 -65
rect 822 -67 824 -65
rect 851 -73 853 -71
rect 813 -80 815 -78
rect 901 -69 903 -67
rect 911 -72 913 -70
rect 921 -80 923 -78
rect 931 -73 933 -71
rect 941 -73 943 -71
rect 931 -80 933 -78
rect 958 -66 960 -64
rect 992 -66 994 -64
rect 1009 -73 1011 -71
rect 1019 -73 1021 -71
rect 1019 -80 1021 -78
rect 1029 -80 1031 -78
rect 1039 -72 1041 -70
rect 1049 -69 1051 -67
rect 1070 -67 1072 -65
rect 1089 -67 1091 -65
rect 1118 -73 1120 -71
rect 1080 -80 1082 -78
rect 1168 -69 1170 -67
rect 1178 -72 1180 -70
rect 1188 -80 1190 -78
rect 1198 -73 1200 -71
rect 1208 -73 1210 -71
rect 1198 -80 1200 -78
rect 1225 -66 1227 -64
rect 1259 -66 1261 -64
rect 1276 -73 1278 -71
rect 1286 -73 1288 -71
rect 1286 -80 1288 -78
rect 1296 -80 1298 -78
rect 1306 -72 1308 -70
rect 1316 -69 1318 -67
rect 1337 -67 1339 -65
rect 1356 -67 1358 -65
rect 1385 -73 1387 -71
rect 1347 -80 1349 -78
rect 1435 -69 1437 -67
rect 1445 -72 1447 -70
rect 1455 -80 1457 -78
rect 1465 -73 1467 -71
rect 1475 -73 1477 -71
rect 1465 -80 1467 -78
rect 1492 -66 1494 -64
rect 1526 -66 1528 -64
rect 1543 -73 1545 -71
rect 1553 -73 1555 -71
rect 1553 -80 1555 -78
rect 1563 -80 1565 -78
rect 1573 -72 1575 -70
rect 1583 -69 1585 -67
rect 1604 -67 1606 -65
rect 1623 -67 1625 -65
rect 1652 -73 1654 -71
rect 1614 -80 1616 -78
rect 1702 -69 1704 -67
rect 1712 -72 1714 -70
rect 1722 -80 1724 -78
rect 1732 -73 1734 -71
rect 1742 -73 1744 -71
rect 1732 -80 1734 -78
rect 1759 -66 1761 -64
rect 1793 -66 1795 -64
rect 1810 -73 1812 -71
rect 1820 -73 1822 -71
rect 1820 -80 1822 -78
rect 1830 -80 1832 -78
rect 1840 -72 1842 -70
rect 1850 -69 1852 -67
rect 1871 -67 1873 -65
rect 1890 -67 1892 -65
rect 1928 -72 1930 -70
rect 1881 -80 1883 -78
rect 1914 -80 1916 -78
rect 1940 -75 1942 -73
rect 1988 -69 1990 -67
rect 1998 -72 2000 -70
rect 2008 -80 2010 -78
rect 2018 -73 2020 -71
rect 2028 -73 2030 -71
rect 2018 -80 2020 -78
rect 2045 -66 2047 -64
rect 2079 -66 2081 -64
rect 2096 -73 2098 -71
rect 2106 -73 2108 -71
rect 2106 -80 2108 -78
rect 2116 -80 2118 -78
rect 2126 -72 2128 -70
rect 2136 -69 2138 -67
rect 2157 -67 2159 -65
rect 2176 -67 2178 -65
rect 2167 -80 2169 -78
rect 2201 -74 2203 -72
rect 2211 -74 2213 -72
rect 2228 -72 2230 -70
rect 2245 -72 2247 -70
rect 2269 -74 2271 -72
rect 2279 -74 2281 -72
rect 2296 -72 2298 -70
rect 2313 -72 2315 -70
rect 10 -185 12 -183
rect 50 -185 52 -183
rect 100 -189 102 -187
rect 110 -186 112 -184
rect 120 -178 122 -176
rect 130 -178 132 -176
rect 130 -185 132 -183
rect 140 -185 142 -183
rect 157 -192 159 -190
rect 191 -192 193 -190
rect 218 -178 220 -176
rect 208 -185 210 -183
rect 218 -185 220 -183
rect 228 -178 230 -176
rect 279 -178 281 -176
rect 238 -186 240 -184
rect 248 -189 250 -187
rect 269 -191 271 -189
rect 317 -185 319 -183
rect 288 -191 290 -189
rect 367 -189 369 -187
rect 377 -186 379 -184
rect 387 -178 389 -176
rect 397 -178 399 -176
rect 397 -185 399 -183
rect 407 -185 409 -183
rect 424 -192 426 -190
rect 458 -192 460 -190
rect 485 -178 487 -176
rect 475 -185 477 -183
rect 485 -185 487 -183
rect 495 -178 497 -176
rect 546 -178 548 -176
rect 505 -186 507 -184
rect 515 -189 517 -187
rect 536 -191 538 -189
rect 584 -185 586 -183
rect 555 -191 557 -189
rect 634 -189 636 -187
rect 644 -186 646 -184
rect 654 -178 656 -176
rect 664 -178 666 -176
rect 664 -185 666 -183
rect 674 -185 676 -183
rect 691 -192 693 -190
rect 725 -192 727 -190
rect 752 -178 754 -176
rect 742 -185 744 -183
rect 752 -185 754 -183
rect 762 -178 764 -176
rect 813 -178 815 -176
rect 772 -186 774 -184
rect 782 -189 784 -187
rect 803 -191 805 -189
rect 851 -185 853 -183
rect 822 -191 824 -189
rect 901 -189 903 -187
rect 911 -186 913 -184
rect 921 -178 923 -176
rect 931 -178 933 -176
rect 931 -185 933 -183
rect 941 -185 943 -183
rect 958 -192 960 -190
rect 992 -192 994 -190
rect 1019 -178 1021 -176
rect 1009 -185 1011 -183
rect 1019 -185 1021 -183
rect 1029 -178 1031 -176
rect 1080 -178 1082 -176
rect 1039 -186 1041 -184
rect 1049 -189 1051 -187
rect 1070 -191 1072 -189
rect 1118 -185 1120 -183
rect 1089 -191 1091 -189
rect 1168 -189 1170 -187
rect 1178 -186 1180 -184
rect 1188 -178 1190 -176
rect 1198 -178 1200 -176
rect 1198 -185 1200 -183
rect 1208 -185 1210 -183
rect 1225 -192 1227 -190
rect 1259 -192 1261 -190
rect 1286 -178 1288 -176
rect 1276 -185 1278 -183
rect 1286 -185 1288 -183
rect 1296 -178 1298 -176
rect 1347 -178 1349 -176
rect 1306 -186 1308 -184
rect 1316 -189 1318 -187
rect 1337 -191 1339 -189
rect 1385 -185 1387 -183
rect 1356 -191 1358 -189
rect 1435 -189 1437 -187
rect 1445 -186 1447 -184
rect 1455 -178 1457 -176
rect 1465 -178 1467 -176
rect 1465 -185 1467 -183
rect 1475 -185 1477 -183
rect 1492 -192 1494 -190
rect 1526 -192 1528 -190
rect 1553 -178 1555 -176
rect 1543 -185 1545 -183
rect 1553 -185 1555 -183
rect 1563 -178 1565 -176
rect 1614 -178 1616 -176
rect 1573 -186 1575 -184
rect 1583 -189 1585 -187
rect 1604 -191 1606 -189
rect 1652 -185 1654 -183
rect 1623 -191 1625 -189
rect 1702 -189 1704 -187
rect 1712 -186 1714 -184
rect 1722 -178 1724 -176
rect 1732 -178 1734 -176
rect 1732 -185 1734 -183
rect 1742 -185 1744 -183
rect 1759 -192 1761 -190
rect 1793 -192 1795 -190
rect 1820 -178 1822 -176
rect 1810 -185 1812 -183
rect 1820 -185 1822 -183
rect 1830 -178 1832 -176
rect 1881 -178 1883 -176
rect 1840 -186 1842 -184
rect 1850 -189 1852 -187
rect 1914 -178 1916 -176
rect 1871 -191 1873 -189
rect 1928 -186 1930 -184
rect 1940 -183 1942 -181
rect 1890 -191 1892 -189
rect 1988 -189 1990 -187
rect 1998 -186 2000 -184
rect 2008 -178 2010 -176
rect 2018 -178 2020 -176
rect 2018 -185 2020 -183
rect 2028 -185 2030 -183
rect 2045 -192 2047 -190
rect 2079 -192 2081 -190
rect 2106 -178 2108 -176
rect 2096 -185 2098 -183
rect 2106 -185 2108 -183
rect 2116 -178 2118 -176
rect 2167 -178 2169 -176
rect 2126 -186 2128 -184
rect 2136 -189 2138 -187
rect 2157 -191 2159 -189
rect 2201 -184 2203 -182
rect 2211 -184 2213 -182
rect 2176 -191 2178 -189
rect 2228 -186 2230 -184
rect 2245 -186 2247 -184
rect 2269 -184 2271 -182
rect 2279 -184 2281 -182
rect 2296 -186 2298 -184
rect 2313 -186 2315 -184
rect 10 -217 12 -215
rect 50 -217 52 -215
rect 100 -213 102 -211
rect 110 -216 112 -214
rect 120 -224 122 -222
rect 130 -217 132 -215
rect 140 -217 142 -215
rect 130 -224 132 -222
rect 157 -210 159 -208
rect 191 -210 193 -208
rect 208 -217 210 -215
rect 218 -217 220 -215
rect 218 -224 220 -222
rect 228 -224 230 -222
rect 238 -216 240 -214
rect 248 -213 250 -211
rect 269 -211 271 -209
rect 288 -211 290 -209
rect 317 -217 319 -215
rect 279 -224 281 -222
rect 367 -213 369 -211
rect 377 -216 379 -214
rect 387 -224 389 -222
rect 397 -217 399 -215
rect 407 -217 409 -215
rect 397 -224 399 -222
rect 424 -210 426 -208
rect 458 -210 460 -208
rect 475 -217 477 -215
rect 485 -217 487 -215
rect 485 -224 487 -222
rect 495 -224 497 -222
rect 505 -216 507 -214
rect 515 -213 517 -211
rect 536 -211 538 -209
rect 555 -211 557 -209
rect 584 -217 586 -215
rect 546 -224 548 -222
rect 634 -213 636 -211
rect 644 -216 646 -214
rect 654 -224 656 -222
rect 664 -217 666 -215
rect 674 -217 676 -215
rect 664 -224 666 -222
rect 691 -210 693 -208
rect 725 -210 727 -208
rect 742 -217 744 -215
rect 752 -217 754 -215
rect 752 -224 754 -222
rect 762 -224 764 -222
rect 772 -216 774 -214
rect 782 -213 784 -211
rect 803 -211 805 -209
rect 822 -211 824 -209
rect 851 -217 853 -215
rect 813 -224 815 -222
rect 901 -213 903 -211
rect 911 -216 913 -214
rect 921 -224 923 -222
rect 931 -217 933 -215
rect 941 -217 943 -215
rect 931 -224 933 -222
rect 958 -210 960 -208
rect 992 -210 994 -208
rect 1009 -217 1011 -215
rect 1019 -217 1021 -215
rect 1019 -224 1021 -222
rect 1029 -224 1031 -222
rect 1039 -216 1041 -214
rect 1049 -213 1051 -211
rect 1070 -211 1072 -209
rect 1089 -211 1091 -209
rect 1118 -217 1120 -215
rect 1080 -224 1082 -222
rect 1168 -213 1170 -211
rect 1178 -216 1180 -214
rect 1188 -224 1190 -222
rect 1198 -217 1200 -215
rect 1208 -217 1210 -215
rect 1198 -224 1200 -222
rect 1225 -210 1227 -208
rect 1259 -210 1261 -208
rect 1276 -217 1278 -215
rect 1286 -217 1288 -215
rect 1286 -224 1288 -222
rect 1296 -224 1298 -222
rect 1306 -216 1308 -214
rect 1316 -213 1318 -211
rect 1337 -211 1339 -209
rect 1356 -211 1358 -209
rect 1385 -217 1387 -215
rect 1347 -224 1349 -222
rect 1435 -213 1437 -211
rect 1445 -216 1447 -214
rect 1455 -224 1457 -222
rect 1465 -217 1467 -215
rect 1475 -217 1477 -215
rect 1465 -224 1467 -222
rect 1492 -210 1494 -208
rect 1526 -210 1528 -208
rect 1543 -217 1545 -215
rect 1553 -217 1555 -215
rect 1553 -224 1555 -222
rect 1563 -224 1565 -222
rect 1573 -216 1575 -214
rect 1583 -213 1585 -211
rect 1604 -211 1606 -209
rect 1623 -211 1625 -209
rect 1652 -217 1654 -215
rect 1614 -224 1616 -222
rect 1702 -213 1704 -211
rect 1712 -216 1714 -214
rect 1722 -224 1724 -222
rect 1732 -217 1734 -215
rect 1742 -217 1744 -215
rect 1732 -224 1734 -222
rect 1759 -210 1761 -208
rect 1793 -210 1795 -208
rect 1810 -217 1812 -215
rect 1820 -217 1822 -215
rect 1820 -224 1822 -222
rect 1830 -224 1832 -222
rect 1840 -216 1842 -214
rect 1850 -213 1852 -211
rect 1871 -211 1873 -209
rect 1890 -211 1892 -209
rect 1928 -216 1930 -214
rect 1881 -224 1883 -222
rect 1914 -224 1916 -222
rect 1940 -219 1942 -217
rect 1988 -213 1990 -211
rect 1998 -216 2000 -214
rect 2008 -224 2010 -222
rect 2018 -217 2020 -215
rect 2028 -217 2030 -215
rect 2018 -224 2020 -222
rect 2045 -210 2047 -208
rect 2079 -210 2081 -208
rect 2096 -217 2098 -215
rect 2106 -217 2108 -215
rect 2106 -224 2108 -222
rect 2116 -224 2118 -222
rect 2126 -216 2128 -214
rect 2136 -213 2138 -211
rect 2157 -211 2159 -209
rect 2176 -211 2178 -209
rect 2167 -224 2169 -222
rect 2201 -218 2203 -216
rect 2211 -218 2213 -216
rect 2228 -216 2230 -214
rect 2245 -216 2247 -214
rect 2269 -218 2271 -216
rect 2279 -218 2281 -216
rect 2296 -216 2298 -214
rect 2313 -216 2315 -214
<< ndifct1 >>
rect 40 249 42 251
rect 80 249 82 251
rect 90 247 92 249
rect 29 237 31 239
rect 69 237 71 239
rect 168 247 170 249
rect 180 247 182 249
rect 258 247 260 249
rect 299 254 301 256
rect 347 249 349 251
rect 357 247 359 249
rect 336 237 338 239
rect 435 247 437 249
rect 447 247 449 249
rect 525 247 527 249
rect 566 254 568 256
rect 614 249 616 251
rect 624 247 626 249
rect 603 237 605 239
rect 702 247 704 249
rect 714 247 716 249
rect 792 247 794 249
rect 833 254 835 256
rect 881 249 883 251
rect 891 247 893 249
rect 870 237 872 239
rect 969 247 971 249
rect 981 247 983 249
rect 1059 247 1061 249
rect 1100 254 1102 256
rect 1148 249 1150 251
rect 1158 247 1160 249
rect 1137 237 1139 239
rect 1236 247 1238 249
rect 1248 247 1250 249
rect 1326 247 1328 249
rect 1367 254 1369 256
rect 1415 249 1417 251
rect 1425 247 1427 249
rect 1404 237 1406 239
rect 1503 247 1505 249
rect 1515 247 1517 249
rect 1593 247 1595 249
rect 1634 254 1636 256
rect 1682 249 1684 251
rect 1692 247 1694 249
rect 1671 237 1673 239
rect 1770 247 1772 249
rect 1782 247 1784 249
rect 1860 247 1862 249
rect 1901 254 1903 256
rect 1950 247 1952 249
rect 1978 247 1980 249
rect 1968 237 1970 239
rect 2056 247 2058 249
rect 2068 247 2070 249
rect 2146 247 2148 249
rect 2187 254 2189 256
rect 2255 249 2257 251
rect 2323 249 2325 251
rect 29 225 31 227
rect 69 225 71 227
rect 40 213 42 215
rect 80 213 82 215
rect 90 215 92 217
rect 168 215 170 217
rect 180 215 182 217
rect 336 225 338 227
rect 258 215 260 217
rect 299 208 301 210
rect 347 213 349 215
rect 357 215 359 217
rect 435 215 437 217
rect 447 215 449 217
rect 603 225 605 227
rect 525 215 527 217
rect 566 208 568 210
rect 614 213 616 215
rect 624 215 626 217
rect 702 215 704 217
rect 714 215 716 217
rect 870 225 872 227
rect 792 215 794 217
rect 833 208 835 210
rect 881 213 883 215
rect 891 215 893 217
rect 969 215 971 217
rect 981 215 983 217
rect 1137 225 1139 227
rect 1059 215 1061 217
rect 1100 208 1102 210
rect 1148 213 1150 215
rect 1158 215 1160 217
rect 1236 215 1238 217
rect 1248 215 1250 217
rect 1404 225 1406 227
rect 1326 215 1328 217
rect 1367 208 1369 210
rect 1415 213 1417 215
rect 1425 215 1427 217
rect 1503 215 1505 217
rect 1515 215 1517 217
rect 1671 225 1673 227
rect 1593 215 1595 217
rect 1634 208 1636 210
rect 1682 213 1684 215
rect 1692 215 1694 217
rect 1770 215 1772 217
rect 1782 215 1784 217
rect 1968 225 1970 227
rect 1860 215 1862 217
rect 1901 208 1903 210
rect 1950 215 1952 217
rect 1978 215 1980 217
rect 2056 215 2058 217
rect 2068 215 2070 217
rect 2146 215 2148 217
rect 2187 208 2189 210
rect 2255 213 2257 215
rect 2323 213 2325 215
rect 40 105 42 107
rect 80 105 82 107
rect 90 103 92 105
rect 29 93 31 95
rect 69 93 71 95
rect 168 103 170 105
rect 180 103 182 105
rect 258 103 260 105
rect 299 110 301 112
rect 347 105 349 107
rect 357 103 359 105
rect 336 93 338 95
rect 435 103 437 105
rect 447 103 449 105
rect 525 103 527 105
rect 566 110 568 112
rect 614 105 616 107
rect 624 103 626 105
rect 603 93 605 95
rect 702 103 704 105
rect 714 103 716 105
rect 792 103 794 105
rect 833 110 835 112
rect 881 105 883 107
rect 891 103 893 105
rect 870 93 872 95
rect 969 103 971 105
rect 981 103 983 105
rect 1059 103 1061 105
rect 1100 110 1102 112
rect 1148 105 1150 107
rect 1158 103 1160 105
rect 1137 93 1139 95
rect 1236 103 1238 105
rect 1248 103 1250 105
rect 1326 103 1328 105
rect 1367 110 1369 112
rect 1415 105 1417 107
rect 1425 103 1427 105
rect 1404 93 1406 95
rect 1503 103 1505 105
rect 1515 103 1517 105
rect 1593 103 1595 105
rect 1634 110 1636 112
rect 1682 105 1684 107
rect 1692 103 1694 105
rect 1671 93 1673 95
rect 1770 103 1772 105
rect 1782 103 1784 105
rect 1860 103 1862 105
rect 1901 110 1903 112
rect 1950 103 1952 105
rect 1978 103 1980 105
rect 1968 93 1970 95
rect 2056 103 2058 105
rect 2068 103 2070 105
rect 2146 103 2148 105
rect 2187 110 2189 112
rect 2255 105 2257 107
rect 2323 105 2325 107
rect 29 81 31 83
rect 69 81 71 83
rect 40 69 42 71
rect 80 69 82 71
rect 90 71 92 73
rect 168 71 170 73
rect 180 71 182 73
rect 336 81 338 83
rect 258 71 260 73
rect 299 64 301 66
rect 347 69 349 71
rect 357 71 359 73
rect 435 71 437 73
rect 447 71 449 73
rect 603 81 605 83
rect 525 71 527 73
rect 566 64 568 66
rect 614 69 616 71
rect 624 71 626 73
rect 702 71 704 73
rect 714 71 716 73
rect 870 81 872 83
rect 792 71 794 73
rect 833 64 835 66
rect 881 69 883 71
rect 891 71 893 73
rect 969 71 971 73
rect 981 71 983 73
rect 1137 81 1139 83
rect 1059 71 1061 73
rect 1100 64 1102 66
rect 1148 69 1150 71
rect 1158 71 1160 73
rect 1236 71 1238 73
rect 1248 71 1250 73
rect 1404 81 1406 83
rect 1326 71 1328 73
rect 1367 64 1369 66
rect 1415 69 1417 71
rect 1425 71 1427 73
rect 1503 71 1505 73
rect 1515 71 1517 73
rect 1671 81 1673 83
rect 1593 71 1595 73
rect 1634 64 1636 66
rect 1682 69 1684 71
rect 1692 71 1694 73
rect 1770 71 1772 73
rect 1782 71 1784 73
rect 1968 81 1970 83
rect 1860 71 1862 73
rect 1901 64 1903 66
rect 1950 71 1952 73
rect 1978 71 1980 73
rect 2056 71 2058 73
rect 2068 71 2070 73
rect 2146 71 2148 73
rect 2187 64 2189 66
rect 2255 69 2257 71
rect 2323 69 2325 71
rect 40 -39 42 -37
rect 80 -39 82 -37
rect 90 -41 92 -39
rect 29 -51 31 -49
rect 69 -51 71 -49
rect 168 -41 170 -39
rect 180 -41 182 -39
rect 258 -41 260 -39
rect 299 -34 301 -32
rect 347 -39 349 -37
rect 357 -41 359 -39
rect 336 -51 338 -49
rect 435 -41 437 -39
rect 447 -41 449 -39
rect 525 -41 527 -39
rect 566 -34 568 -32
rect 614 -39 616 -37
rect 624 -41 626 -39
rect 603 -51 605 -49
rect 702 -41 704 -39
rect 714 -41 716 -39
rect 792 -41 794 -39
rect 833 -34 835 -32
rect 881 -39 883 -37
rect 891 -41 893 -39
rect 870 -51 872 -49
rect 969 -41 971 -39
rect 981 -41 983 -39
rect 1059 -41 1061 -39
rect 1100 -34 1102 -32
rect 1148 -39 1150 -37
rect 1158 -41 1160 -39
rect 1137 -51 1139 -49
rect 1236 -41 1238 -39
rect 1248 -41 1250 -39
rect 1326 -41 1328 -39
rect 1367 -34 1369 -32
rect 1415 -39 1417 -37
rect 1425 -41 1427 -39
rect 1404 -51 1406 -49
rect 1503 -41 1505 -39
rect 1515 -41 1517 -39
rect 1593 -41 1595 -39
rect 1634 -34 1636 -32
rect 1682 -39 1684 -37
rect 1692 -41 1694 -39
rect 1671 -51 1673 -49
rect 1770 -41 1772 -39
rect 1782 -41 1784 -39
rect 1860 -41 1862 -39
rect 1901 -34 1903 -32
rect 1950 -41 1952 -39
rect 1978 -41 1980 -39
rect 1968 -51 1970 -49
rect 2056 -41 2058 -39
rect 2068 -41 2070 -39
rect 2146 -41 2148 -39
rect 2187 -34 2189 -32
rect 2255 -39 2257 -37
rect 2323 -39 2325 -37
rect 29 -63 31 -61
rect 69 -63 71 -61
rect 40 -75 42 -73
rect 80 -75 82 -73
rect 90 -73 92 -71
rect 168 -73 170 -71
rect 180 -73 182 -71
rect 336 -63 338 -61
rect 258 -73 260 -71
rect 299 -80 301 -78
rect 347 -75 349 -73
rect 357 -73 359 -71
rect 435 -73 437 -71
rect 447 -73 449 -71
rect 603 -63 605 -61
rect 525 -73 527 -71
rect 566 -80 568 -78
rect 614 -75 616 -73
rect 624 -73 626 -71
rect 702 -73 704 -71
rect 714 -73 716 -71
rect 870 -63 872 -61
rect 792 -73 794 -71
rect 833 -80 835 -78
rect 881 -75 883 -73
rect 891 -73 893 -71
rect 969 -73 971 -71
rect 981 -73 983 -71
rect 1137 -63 1139 -61
rect 1059 -73 1061 -71
rect 1100 -80 1102 -78
rect 1148 -75 1150 -73
rect 1158 -73 1160 -71
rect 1236 -73 1238 -71
rect 1248 -73 1250 -71
rect 1404 -63 1406 -61
rect 1326 -73 1328 -71
rect 1367 -80 1369 -78
rect 1415 -75 1417 -73
rect 1425 -73 1427 -71
rect 1503 -73 1505 -71
rect 1515 -73 1517 -71
rect 1671 -63 1673 -61
rect 1593 -73 1595 -71
rect 1634 -80 1636 -78
rect 1682 -75 1684 -73
rect 1692 -73 1694 -71
rect 1770 -73 1772 -71
rect 1782 -73 1784 -71
rect 1968 -63 1970 -61
rect 1860 -73 1862 -71
rect 1901 -80 1903 -78
rect 1950 -73 1952 -71
rect 1978 -73 1980 -71
rect 2056 -73 2058 -71
rect 2068 -73 2070 -71
rect 2146 -73 2148 -71
rect 2187 -80 2189 -78
rect 2255 -75 2257 -73
rect 2323 -75 2325 -73
rect 40 -183 42 -181
rect 80 -183 82 -181
rect 90 -185 92 -183
rect 29 -195 31 -193
rect 69 -195 71 -193
rect 168 -185 170 -183
rect 180 -185 182 -183
rect 258 -185 260 -183
rect 299 -178 301 -176
rect 347 -183 349 -181
rect 357 -185 359 -183
rect 336 -195 338 -193
rect 435 -185 437 -183
rect 447 -185 449 -183
rect 525 -185 527 -183
rect 566 -178 568 -176
rect 614 -183 616 -181
rect 624 -185 626 -183
rect 603 -195 605 -193
rect 702 -185 704 -183
rect 714 -185 716 -183
rect 792 -185 794 -183
rect 833 -178 835 -176
rect 881 -183 883 -181
rect 891 -185 893 -183
rect 870 -195 872 -193
rect 969 -185 971 -183
rect 981 -185 983 -183
rect 1059 -185 1061 -183
rect 1100 -178 1102 -176
rect 1148 -183 1150 -181
rect 1158 -185 1160 -183
rect 1137 -195 1139 -193
rect 1236 -185 1238 -183
rect 1248 -185 1250 -183
rect 1326 -185 1328 -183
rect 1367 -178 1369 -176
rect 1415 -183 1417 -181
rect 1425 -185 1427 -183
rect 1404 -195 1406 -193
rect 1503 -185 1505 -183
rect 1515 -185 1517 -183
rect 1593 -185 1595 -183
rect 1634 -178 1636 -176
rect 1682 -183 1684 -181
rect 1692 -185 1694 -183
rect 1671 -195 1673 -193
rect 1770 -185 1772 -183
rect 1782 -185 1784 -183
rect 1860 -185 1862 -183
rect 1901 -178 1903 -176
rect 1950 -185 1952 -183
rect 1978 -185 1980 -183
rect 1968 -195 1970 -193
rect 2056 -185 2058 -183
rect 2068 -185 2070 -183
rect 2146 -185 2148 -183
rect 2187 -178 2189 -176
rect 2255 -183 2257 -181
rect 2323 -183 2325 -181
rect 29 -207 31 -205
rect 69 -207 71 -205
rect 40 -219 42 -217
rect 80 -219 82 -217
rect 90 -217 92 -215
rect 168 -217 170 -215
rect 180 -217 182 -215
rect 336 -207 338 -205
rect 258 -217 260 -215
rect 299 -224 301 -222
rect 347 -219 349 -217
rect 357 -217 359 -215
rect 435 -217 437 -215
rect 447 -217 449 -215
rect 603 -207 605 -205
rect 525 -217 527 -215
rect 566 -224 568 -222
rect 614 -219 616 -217
rect 624 -217 626 -215
rect 702 -217 704 -215
rect 714 -217 716 -215
rect 870 -207 872 -205
rect 792 -217 794 -215
rect 833 -224 835 -222
rect 881 -219 883 -217
rect 891 -217 893 -215
rect 969 -217 971 -215
rect 981 -217 983 -215
rect 1137 -207 1139 -205
rect 1059 -217 1061 -215
rect 1100 -224 1102 -222
rect 1148 -219 1150 -217
rect 1158 -217 1160 -215
rect 1236 -217 1238 -215
rect 1248 -217 1250 -215
rect 1404 -207 1406 -205
rect 1326 -217 1328 -215
rect 1367 -224 1369 -222
rect 1415 -219 1417 -217
rect 1425 -217 1427 -215
rect 1503 -217 1505 -215
rect 1515 -217 1517 -215
rect 1671 -207 1673 -205
rect 1593 -217 1595 -215
rect 1634 -224 1636 -222
rect 1682 -219 1684 -217
rect 1692 -217 1694 -215
rect 1770 -217 1772 -215
rect 1782 -217 1784 -215
rect 1968 -207 1970 -205
rect 1860 -217 1862 -215
rect 1901 -224 1903 -222
rect 1950 -217 1952 -215
rect 1978 -217 1980 -215
rect 2056 -217 2058 -215
rect 2068 -217 2070 -215
rect 2146 -217 2148 -215
rect 2187 -224 2189 -222
rect 2255 -219 2257 -217
rect 2323 -219 2325 -217
<< ntiect1 >>
rect 39 297 41 299
rect 79 297 81 299
rect 298 297 300 299
rect 346 297 348 299
rect 565 297 567 299
rect 613 297 615 299
rect 832 297 834 299
rect 880 297 882 299
rect 1099 297 1101 299
rect 1147 297 1149 299
rect 1366 297 1368 299
rect 1414 297 1416 299
rect 1633 297 1635 299
rect 1681 297 1683 299
rect 1900 297 1902 299
rect 1948 297 1950 299
rect 2186 297 2188 299
rect 39 165 41 167
rect 79 165 81 167
rect 298 165 300 167
rect 346 165 348 167
rect 565 165 567 167
rect 613 165 615 167
rect 832 165 834 167
rect 880 165 882 167
rect 1099 165 1101 167
rect 1147 165 1149 167
rect 1366 165 1368 167
rect 1414 165 1416 167
rect 1633 165 1635 167
rect 1681 165 1683 167
rect 1900 165 1902 167
rect 1948 165 1950 167
rect 2186 165 2188 167
rect 39 153 41 155
rect 79 153 81 155
rect 298 153 300 155
rect 346 153 348 155
rect 565 153 567 155
rect 613 153 615 155
rect 832 153 834 155
rect 880 153 882 155
rect 1099 153 1101 155
rect 1147 153 1149 155
rect 1366 153 1368 155
rect 1414 153 1416 155
rect 1633 153 1635 155
rect 1681 153 1683 155
rect 1900 153 1902 155
rect 1948 153 1950 155
rect 2186 153 2188 155
rect 39 21 41 23
rect 79 21 81 23
rect 298 21 300 23
rect 346 21 348 23
rect 565 21 567 23
rect 613 21 615 23
rect 832 21 834 23
rect 880 21 882 23
rect 1099 21 1101 23
rect 1147 21 1149 23
rect 1366 21 1368 23
rect 1414 21 1416 23
rect 1633 21 1635 23
rect 1681 21 1683 23
rect 1900 21 1902 23
rect 1948 21 1950 23
rect 2186 21 2188 23
rect 39 9 41 11
rect 79 9 81 11
rect 298 9 300 11
rect 346 9 348 11
rect 565 9 567 11
rect 613 9 615 11
rect 832 9 834 11
rect 880 9 882 11
rect 1099 9 1101 11
rect 1147 9 1149 11
rect 1366 9 1368 11
rect 1414 9 1416 11
rect 1633 9 1635 11
rect 1681 9 1683 11
rect 1900 9 1902 11
rect 1948 9 1950 11
rect 2186 9 2188 11
rect 39 -123 41 -121
rect 79 -123 81 -121
rect 298 -123 300 -121
rect 346 -123 348 -121
rect 565 -123 567 -121
rect 613 -123 615 -121
rect 832 -123 834 -121
rect 880 -123 882 -121
rect 1099 -123 1101 -121
rect 1147 -123 1149 -121
rect 1366 -123 1368 -121
rect 1414 -123 1416 -121
rect 1633 -123 1635 -121
rect 1681 -123 1683 -121
rect 1900 -123 1902 -121
rect 1948 -123 1950 -121
rect 2186 -123 2188 -121
rect 39 -135 41 -133
rect 79 -135 81 -133
rect 298 -135 300 -133
rect 346 -135 348 -133
rect 565 -135 567 -133
rect 613 -135 615 -133
rect 832 -135 834 -133
rect 880 -135 882 -133
rect 1099 -135 1101 -133
rect 1147 -135 1149 -133
rect 1366 -135 1368 -133
rect 1414 -135 1416 -133
rect 1633 -135 1635 -133
rect 1681 -135 1683 -133
rect 1900 -135 1902 -133
rect 1948 -135 1950 -133
rect 2186 -135 2188 -133
rect 39 -267 41 -265
rect 79 -267 81 -265
rect 298 -267 300 -265
rect 346 -267 348 -265
rect 565 -267 567 -265
rect 613 -267 615 -265
rect 832 -267 834 -265
rect 880 -267 882 -265
rect 1099 -267 1101 -265
rect 1147 -267 1149 -265
rect 1366 -267 1368 -265
rect 1414 -267 1416 -265
rect 1633 -267 1635 -265
rect 1681 -267 1683 -265
rect 1900 -267 1902 -265
rect 1948 -267 1950 -265
rect 2186 -267 2188 -265
<< ptiect1 >>
rect 39 237 41 239
rect 79 237 81 239
rect 298 237 300 239
rect 346 237 348 239
rect 565 237 567 239
rect 613 237 615 239
rect 832 237 834 239
rect 880 237 882 239
rect 1099 237 1101 239
rect 1147 237 1149 239
rect 1366 237 1368 239
rect 1414 237 1416 239
rect 1633 237 1635 239
rect 1681 237 1683 239
rect 1900 237 1902 239
rect 1915 237 1917 239
rect 2186 237 2188 239
rect 39 225 41 227
rect 79 225 81 227
rect 298 225 300 227
rect 346 225 348 227
rect 565 225 567 227
rect 613 225 615 227
rect 832 225 834 227
rect 880 225 882 227
rect 1099 225 1101 227
rect 1147 225 1149 227
rect 1366 225 1368 227
rect 1414 225 1416 227
rect 1633 225 1635 227
rect 1681 225 1683 227
rect 1900 225 1902 227
rect 1915 225 1917 227
rect 2186 225 2188 227
rect 39 93 41 95
rect 79 93 81 95
rect 298 93 300 95
rect 346 93 348 95
rect 565 93 567 95
rect 613 93 615 95
rect 832 93 834 95
rect 880 93 882 95
rect 1099 93 1101 95
rect 1147 93 1149 95
rect 1366 93 1368 95
rect 1414 93 1416 95
rect 1633 93 1635 95
rect 1681 93 1683 95
rect 1900 93 1902 95
rect 1915 93 1917 95
rect 2186 93 2188 95
rect 39 81 41 83
rect 79 81 81 83
rect 298 81 300 83
rect 346 81 348 83
rect 565 81 567 83
rect 613 81 615 83
rect 832 81 834 83
rect 880 81 882 83
rect 1099 81 1101 83
rect 1147 81 1149 83
rect 1366 81 1368 83
rect 1414 81 1416 83
rect 1633 81 1635 83
rect 1681 81 1683 83
rect 1900 81 1902 83
rect 1915 81 1917 83
rect 2186 81 2188 83
rect 39 -51 41 -49
rect 79 -51 81 -49
rect 298 -51 300 -49
rect 346 -51 348 -49
rect 565 -51 567 -49
rect 613 -51 615 -49
rect 832 -51 834 -49
rect 880 -51 882 -49
rect 1099 -51 1101 -49
rect 1147 -51 1149 -49
rect 1366 -51 1368 -49
rect 1414 -51 1416 -49
rect 1633 -51 1635 -49
rect 1681 -51 1683 -49
rect 1900 -51 1902 -49
rect 1915 -51 1917 -49
rect 2186 -51 2188 -49
rect 39 -63 41 -61
rect 79 -63 81 -61
rect 298 -63 300 -61
rect 346 -63 348 -61
rect 565 -63 567 -61
rect 613 -63 615 -61
rect 832 -63 834 -61
rect 880 -63 882 -61
rect 1099 -63 1101 -61
rect 1147 -63 1149 -61
rect 1366 -63 1368 -61
rect 1414 -63 1416 -61
rect 1633 -63 1635 -61
rect 1681 -63 1683 -61
rect 1900 -63 1902 -61
rect 1915 -63 1917 -61
rect 2186 -63 2188 -61
rect 39 -195 41 -193
rect 79 -195 81 -193
rect 298 -195 300 -193
rect 346 -195 348 -193
rect 565 -195 567 -193
rect 613 -195 615 -193
rect 832 -195 834 -193
rect 880 -195 882 -193
rect 1099 -195 1101 -193
rect 1147 -195 1149 -193
rect 1366 -195 1368 -193
rect 1414 -195 1416 -193
rect 1633 -195 1635 -193
rect 1681 -195 1683 -193
rect 1900 -195 1902 -193
rect 1915 -195 1917 -193
rect 2186 -195 2188 -193
rect 39 -207 41 -205
rect 79 -207 81 -205
rect 298 -207 300 -205
rect 346 -207 348 -205
rect 565 -207 567 -205
rect 613 -207 615 -205
rect 832 -207 834 -205
rect 880 -207 882 -205
rect 1099 -207 1101 -205
rect 1147 -207 1149 -205
rect 1366 -207 1368 -205
rect 1414 -207 1416 -205
rect 1633 -207 1635 -205
rect 1681 -207 1683 -205
rect 1900 -207 1902 -205
rect 1915 -207 1917 -205
rect 2186 -207 2188 -205
<< pdifct0 >>
rect 10 287 12 289
rect 20 287 22 289
rect 20 280 22 282
rect 30 285 32 287
rect 50 287 52 289
rect 60 287 62 289
rect 60 280 62 282
rect 70 285 72 287
rect 101 294 103 296
rect 113 275 115 277
rect 136 294 138 296
rect 136 287 138 289
rect 148 286 150 288
rect 148 279 150 281
rect 158 294 160 296
rect 158 287 160 289
rect 190 294 192 296
rect 190 287 192 289
rect 200 286 202 288
rect 200 279 202 281
rect 212 294 214 296
rect 212 287 214 289
rect 247 294 249 296
rect 235 275 237 277
rect 269 287 271 289
rect 288 294 290 296
rect 317 287 319 289
rect 327 287 329 289
rect 327 280 329 282
rect 337 285 339 287
rect 368 294 370 296
rect 380 275 382 277
rect 403 294 405 296
rect 403 287 405 289
rect 415 286 417 288
rect 415 279 417 281
rect 425 294 427 296
rect 425 287 427 289
rect 457 294 459 296
rect 457 287 459 289
rect 467 286 469 288
rect 467 279 469 281
rect 479 294 481 296
rect 479 287 481 289
rect 514 294 516 296
rect 502 275 504 277
rect 536 287 538 289
rect 555 294 557 296
rect 584 287 586 289
rect 594 287 596 289
rect 594 280 596 282
rect 604 285 606 287
rect 635 294 637 296
rect 647 275 649 277
rect 670 294 672 296
rect 670 287 672 289
rect 682 286 684 288
rect 682 279 684 281
rect 692 294 694 296
rect 692 287 694 289
rect 724 294 726 296
rect 724 287 726 289
rect 734 286 736 288
rect 734 279 736 281
rect 746 294 748 296
rect 746 287 748 289
rect 781 294 783 296
rect 769 275 771 277
rect 803 287 805 289
rect 822 294 824 296
rect 851 287 853 289
rect 861 287 863 289
rect 861 280 863 282
rect 871 285 873 287
rect 902 294 904 296
rect 914 275 916 277
rect 937 294 939 296
rect 937 287 939 289
rect 949 286 951 288
rect 949 279 951 281
rect 959 294 961 296
rect 959 287 961 289
rect 991 294 993 296
rect 991 287 993 289
rect 1001 286 1003 288
rect 1001 279 1003 281
rect 1013 294 1015 296
rect 1013 287 1015 289
rect 1048 294 1050 296
rect 1036 275 1038 277
rect 1070 287 1072 289
rect 1089 294 1091 296
rect 1118 287 1120 289
rect 1128 287 1130 289
rect 1128 280 1130 282
rect 1138 285 1140 287
rect 1169 294 1171 296
rect 1181 275 1183 277
rect 1204 294 1206 296
rect 1204 287 1206 289
rect 1216 286 1218 288
rect 1216 279 1218 281
rect 1226 294 1228 296
rect 1226 287 1228 289
rect 1258 294 1260 296
rect 1258 287 1260 289
rect 1268 286 1270 288
rect 1268 279 1270 281
rect 1280 294 1282 296
rect 1280 287 1282 289
rect 1315 294 1317 296
rect 1303 275 1305 277
rect 1337 287 1339 289
rect 1356 294 1358 296
rect 1385 287 1387 289
rect 1395 287 1397 289
rect 1395 280 1397 282
rect 1405 285 1407 287
rect 1436 294 1438 296
rect 1448 275 1450 277
rect 1471 294 1473 296
rect 1471 287 1473 289
rect 1483 286 1485 288
rect 1483 279 1485 281
rect 1493 294 1495 296
rect 1493 287 1495 289
rect 1525 294 1527 296
rect 1525 287 1527 289
rect 1535 286 1537 288
rect 1535 279 1537 281
rect 1547 294 1549 296
rect 1547 287 1549 289
rect 1582 294 1584 296
rect 1570 275 1572 277
rect 1604 287 1606 289
rect 1623 294 1625 296
rect 1652 287 1654 289
rect 1662 287 1664 289
rect 1662 280 1664 282
rect 1672 285 1674 287
rect 1703 294 1705 296
rect 1715 275 1717 277
rect 1738 294 1740 296
rect 1738 287 1740 289
rect 1750 286 1752 288
rect 1750 279 1752 281
rect 1760 294 1762 296
rect 1760 287 1762 289
rect 1792 294 1794 296
rect 1792 287 1794 289
rect 1802 286 1804 288
rect 1802 279 1804 281
rect 1814 294 1816 296
rect 1814 287 1816 289
rect 1849 294 1851 296
rect 1837 275 1839 277
rect 1871 287 1873 289
rect 1890 294 1892 296
rect 1922 273 1924 275
rect 1932 294 1934 296
rect 1932 287 1934 289
rect 1948 280 1950 282
rect 1948 273 1950 275
rect 1968 288 1970 290
rect 1989 294 1991 296
rect 2001 275 2003 277
rect 2024 294 2026 296
rect 2024 287 2026 289
rect 2036 286 2038 288
rect 2036 279 2038 281
rect 2046 294 2048 296
rect 2046 287 2048 289
rect 2078 294 2080 296
rect 2078 287 2080 289
rect 2088 286 2090 288
rect 2088 279 2090 281
rect 2100 294 2102 296
rect 2100 287 2102 289
rect 2135 294 2137 296
rect 2123 275 2125 277
rect 2157 287 2159 289
rect 2176 294 2178 296
rect 2211 294 2213 296
rect 2228 284 2230 286
rect 2245 294 2247 296
rect 2201 272 2203 274
rect 2279 294 2281 296
rect 2296 284 2298 286
rect 2313 294 2315 296
rect 2269 272 2271 274
rect 10 175 12 177
rect 20 182 22 184
rect 20 175 22 177
rect 30 177 32 179
rect 50 175 52 177
rect 60 182 62 184
rect 60 175 62 177
rect 70 177 72 179
rect 113 187 115 189
rect 101 168 103 170
rect 136 175 138 177
rect 136 168 138 170
rect 148 183 150 185
rect 148 176 150 178
rect 158 175 160 177
rect 158 168 160 170
rect 190 175 192 177
rect 190 168 192 170
rect 200 183 202 185
rect 200 176 202 178
rect 212 175 214 177
rect 212 168 214 170
rect 235 187 237 189
rect 247 168 249 170
rect 269 175 271 177
rect 317 175 319 177
rect 327 182 329 184
rect 327 175 329 177
rect 337 177 339 179
rect 288 168 290 170
rect 380 187 382 189
rect 368 168 370 170
rect 403 175 405 177
rect 403 168 405 170
rect 415 183 417 185
rect 415 176 417 178
rect 425 175 427 177
rect 425 168 427 170
rect 457 175 459 177
rect 457 168 459 170
rect 467 183 469 185
rect 467 176 469 178
rect 479 175 481 177
rect 479 168 481 170
rect 502 187 504 189
rect 514 168 516 170
rect 536 175 538 177
rect 584 175 586 177
rect 594 182 596 184
rect 594 175 596 177
rect 604 177 606 179
rect 555 168 557 170
rect 647 187 649 189
rect 635 168 637 170
rect 670 175 672 177
rect 670 168 672 170
rect 682 183 684 185
rect 682 176 684 178
rect 692 175 694 177
rect 692 168 694 170
rect 724 175 726 177
rect 724 168 726 170
rect 734 183 736 185
rect 734 176 736 178
rect 746 175 748 177
rect 746 168 748 170
rect 769 187 771 189
rect 781 168 783 170
rect 803 175 805 177
rect 851 175 853 177
rect 861 182 863 184
rect 861 175 863 177
rect 871 177 873 179
rect 822 168 824 170
rect 914 187 916 189
rect 902 168 904 170
rect 937 175 939 177
rect 937 168 939 170
rect 949 183 951 185
rect 949 176 951 178
rect 959 175 961 177
rect 959 168 961 170
rect 991 175 993 177
rect 991 168 993 170
rect 1001 183 1003 185
rect 1001 176 1003 178
rect 1013 175 1015 177
rect 1013 168 1015 170
rect 1036 187 1038 189
rect 1048 168 1050 170
rect 1070 175 1072 177
rect 1118 175 1120 177
rect 1128 182 1130 184
rect 1128 175 1130 177
rect 1138 177 1140 179
rect 1089 168 1091 170
rect 1181 187 1183 189
rect 1169 168 1171 170
rect 1204 175 1206 177
rect 1204 168 1206 170
rect 1216 183 1218 185
rect 1216 176 1218 178
rect 1226 175 1228 177
rect 1226 168 1228 170
rect 1258 175 1260 177
rect 1258 168 1260 170
rect 1268 183 1270 185
rect 1268 176 1270 178
rect 1280 175 1282 177
rect 1280 168 1282 170
rect 1303 187 1305 189
rect 1315 168 1317 170
rect 1337 175 1339 177
rect 1385 175 1387 177
rect 1395 182 1397 184
rect 1395 175 1397 177
rect 1405 177 1407 179
rect 1356 168 1358 170
rect 1448 187 1450 189
rect 1436 168 1438 170
rect 1471 175 1473 177
rect 1471 168 1473 170
rect 1483 183 1485 185
rect 1483 176 1485 178
rect 1493 175 1495 177
rect 1493 168 1495 170
rect 1525 175 1527 177
rect 1525 168 1527 170
rect 1535 183 1537 185
rect 1535 176 1537 178
rect 1547 175 1549 177
rect 1547 168 1549 170
rect 1570 187 1572 189
rect 1582 168 1584 170
rect 1604 175 1606 177
rect 1652 175 1654 177
rect 1662 182 1664 184
rect 1662 175 1664 177
rect 1672 177 1674 179
rect 1623 168 1625 170
rect 1715 187 1717 189
rect 1703 168 1705 170
rect 1738 175 1740 177
rect 1738 168 1740 170
rect 1750 183 1752 185
rect 1750 176 1752 178
rect 1760 175 1762 177
rect 1760 168 1762 170
rect 1792 175 1794 177
rect 1792 168 1794 170
rect 1802 183 1804 185
rect 1802 176 1804 178
rect 1814 175 1816 177
rect 1814 168 1816 170
rect 1837 187 1839 189
rect 1849 168 1851 170
rect 1871 175 1873 177
rect 1922 189 1924 191
rect 1890 168 1892 170
rect 1932 175 1934 177
rect 1948 189 1950 191
rect 1948 182 1950 184
rect 1932 168 1934 170
rect 1968 174 1970 176
rect 2001 187 2003 189
rect 1989 168 1991 170
rect 2024 175 2026 177
rect 2024 168 2026 170
rect 2036 183 2038 185
rect 2036 176 2038 178
rect 2046 175 2048 177
rect 2046 168 2048 170
rect 2078 175 2080 177
rect 2078 168 2080 170
rect 2088 183 2090 185
rect 2088 176 2090 178
rect 2100 175 2102 177
rect 2100 168 2102 170
rect 2123 187 2125 189
rect 2135 168 2137 170
rect 2157 175 2159 177
rect 2201 190 2203 192
rect 2269 190 2271 192
rect 2176 168 2178 170
rect 2211 168 2213 170
rect 2228 178 2230 180
rect 2245 168 2247 170
rect 2279 168 2281 170
rect 2296 178 2298 180
rect 2313 168 2315 170
rect 10 143 12 145
rect 20 143 22 145
rect 20 136 22 138
rect 30 141 32 143
rect 50 143 52 145
rect 60 143 62 145
rect 60 136 62 138
rect 70 141 72 143
rect 101 150 103 152
rect 113 131 115 133
rect 136 150 138 152
rect 136 143 138 145
rect 148 142 150 144
rect 148 135 150 137
rect 158 150 160 152
rect 158 143 160 145
rect 190 150 192 152
rect 190 143 192 145
rect 200 142 202 144
rect 200 135 202 137
rect 212 150 214 152
rect 212 143 214 145
rect 247 150 249 152
rect 235 131 237 133
rect 269 143 271 145
rect 288 150 290 152
rect 317 143 319 145
rect 327 143 329 145
rect 327 136 329 138
rect 337 141 339 143
rect 368 150 370 152
rect 380 131 382 133
rect 403 150 405 152
rect 403 143 405 145
rect 415 142 417 144
rect 415 135 417 137
rect 425 150 427 152
rect 425 143 427 145
rect 457 150 459 152
rect 457 143 459 145
rect 467 142 469 144
rect 467 135 469 137
rect 479 150 481 152
rect 479 143 481 145
rect 514 150 516 152
rect 502 131 504 133
rect 536 143 538 145
rect 555 150 557 152
rect 584 143 586 145
rect 594 143 596 145
rect 594 136 596 138
rect 604 141 606 143
rect 635 150 637 152
rect 647 131 649 133
rect 670 150 672 152
rect 670 143 672 145
rect 682 142 684 144
rect 682 135 684 137
rect 692 150 694 152
rect 692 143 694 145
rect 724 150 726 152
rect 724 143 726 145
rect 734 142 736 144
rect 734 135 736 137
rect 746 150 748 152
rect 746 143 748 145
rect 781 150 783 152
rect 769 131 771 133
rect 803 143 805 145
rect 822 150 824 152
rect 851 143 853 145
rect 861 143 863 145
rect 861 136 863 138
rect 871 141 873 143
rect 902 150 904 152
rect 914 131 916 133
rect 937 150 939 152
rect 937 143 939 145
rect 949 142 951 144
rect 949 135 951 137
rect 959 150 961 152
rect 959 143 961 145
rect 991 150 993 152
rect 991 143 993 145
rect 1001 142 1003 144
rect 1001 135 1003 137
rect 1013 150 1015 152
rect 1013 143 1015 145
rect 1048 150 1050 152
rect 1036 131 1038 133
rect 1070 143 1072 145
rect 1089 150 1091 152
rect 1118 143 1120 145
rect 1128 143 1130 145
rect 1128 136 1130 138
rect 1138 141 1140 143
rect 1169 150 1171 152
rect 1181 131 1183 133
rect 1204 150 1206 152
rect 1204 143 1206 145
rect 1216 142 1218 144
rect 1216 135 1218 137
rect 1226 150 1228 152
rect 1226 143 1228 145
rect 1258 150 1260 152
rect 1258 143 1260 145
rect 1268 142 1270 144
rect 1268 135 1270 137
rect 1280 150 1282 152
rect 1280 143 1282 145
rect 1315 150 1317 152
rect 1303 131 1305 133
rect 1337 143 1339 145
rect 1356 150 1358 152
rect 1385 143 1387 145
rect 1395 143 1397 145
rect 1395 136 1397 138
rect 1405 141 1407 143
rect 1436 150 1438 152
rect 1448 131 1450 133
rect 1471 150 1473 152
rect 1471 143 1473 145
rect 1483 142 1485 144
rect 1483 135 1485 137
rect 1493 150 1495 152
rect 1493 143 1495 145
rect 1525 150 1527 152
rect 1525 143 1527 145
rect 1535 142 1537 144
rect 1535 135 1537 137
rect 1547 150 1549 152
rect 1547 143 1549 145
rect 1582 150 1584 152
rect 1570 131 1572 133
rect 1604 143 1606 145
rect 1623 150 1625 152
rect 1652 143 1654 145
rect 1662 143 1664 145
rect 1662 136 1664 138
rect 1672 141 1674 143
rect 1703 150 1705 152
rect 1715 131 1717 133
rect 1738 150 1740 152
rect 1738 143 1740 145
rect 1750 142 1752 144
rect 1750 135 1752 137
rect 1760 150 1762 152
rect 1760 143 1762 145
rect 1792 150 1794 152
rect 1792 143 1794 145
rect 1802 142 1804 144
rect 1802 135 1804 137
rect 1814 150 1816 152
rect 1814 143 1816 145
rect 1849 150 1851 152
rect 1837 131 1839 133
rect 1871 143 1873 145
rect 1890 150 1892 152
rect 1922 129 1924 131
rect 1932 150 1934 152
rect 1932 143 1934 145
rect 1948 136 1950 138
rect 1948 129 1950 131
rect 1968 144 1970 146
rect 1989 150 1991 152
rect 2001 131 2003 133
rect 2024 150 2026 152
rect 2024 143 2026 145
rect 2036 142 2038 144
rect 2036 135 2038 137
rect 2046 150 2048 152
rect 2046 143 2048 145
rect 2078 150 2080 152
rect 2078 143 2080 145
rect 2088 142 2090 144
rect 2088 135 2090 137
rect 2100 150 2102 152
rect 2100 143 2102 145
rect 2135 150 2137 152
rect 2123 131 2125 133
rect 2157 143 2159 145
rect 2176 150 2178 152
rect 2211 150 2213 152
rect 2228 140 2230 142
rect 2245 150 2247 152
rect 2201 128 2203 130
rect 2279 150 2281 152
rect 2296 140 2298 142
rect 2313 150 2315 152
rect 2269 128 2271 130
rect 10 31 12 33
rect 20 38 22 40
rect 20 31 22 33
rect 30 33 32 35
rect 50 31 52 33
rect 60 38 62 40
rect 60 31 62 33
rect 70 33 72 35
rect 113 43 115 45
rect 101 24 103 26
rect 136 31 138 33
rect 136 24 138 26
rect 148 39 150 41
rect 148 32 150 34
rect 158 31 160 33
rect 158 24 160 26
rect 190 31 192 33
rect 190 24 192 26
rect 200 39 202 41
rect 200 32 202 34
rect 212 31 214 33
rect 212 24 214 26
rect 235 43 237 45
rect 247 24 249 26
rect 269 31 271 33
rect 317 31 319 33
rect 327 38 329 40
rect 327 31 329 33
rect 337 33 339 35
rect 288 24 290 26
rect 380 43 382 45
rect 368 24 370 26
rect 403 31 405 33
rect 403 24 405 26
rect 415 39 417 41
rect 415 32 417 34
rect 425 31 427 33
rect 425 24 427 26
rect 457 31 459 33
rect 457 24 459 26
rect 467 39 469 41
rect 467 32 469 34
rect 479 31 481 33
rect 479 24 481 26
rect 502 43 504 45
rect 514 24 516 26
rect 536 31 538 33
rect 584 31 586 33
rect 594 38 596 40
rect 594 31 596 33
rect 604 33 606 35
rect 555 24 557 26
rect 647 43 649 45
rect 635 24 637 26
rect 670 31 672 33
rect 670 24 672 26
rect 682 39 684 41
rect 682 32 684 34
rect 692 31 694 33
rect 692 24 694 26
rect 724 31 726 33
rect 724 24 726 26
rect 734 39 736 41
rect 734 32 736 34
rect 746 31 748 33
rect 746 24 748 26
rect 769 43 771 45
rect 781 24 783 26
rect 803 31 805 33
rect 851 31 853 33
rect 861 38 863 40
rect 861 31 863 33
rect 871 33 873 35
rect 822 24 824 26
rect 914 43 916 45
rect 902 24 904 26
rect 937 31 939 33
rect 937 24 939 26
rect 949 39 951 41
rect 949 32 951 34
rect 959 31 961 33
rect 959 24 961 26
rect 991 31 993 33
rect 991 24 993 26
rect 1001 39 1003 41
rect 1001 32 1003 34
rect 1013 31 1015 33
rect 1013 24 1015 26
rect 1036 43 1038 45
rect 1048 24 1050 26
rect 1070 31 1072 33
rect 1118 31 1120 33
rect 1128 38 1130 40
rect 1128 31 1130 33
rect 1138 33 1140 35
rect 1089 24 1091 26
rect 1181 43 1183 45
rect 1169 24 1171 26
rect 1204 31 1206 33
rect 1204 24 1206 26
rect 1216 39 1218 41
rect 1216 32 1218 34
rect 1226 31 1228 33
rect 1226 24 1228 26
rect 1258 31 1260 33
rect 1258 24 1260 26
rect 1268 39 1270 41
rect 1268 32 1270 34
rect 1280 31 1282 33
rect 1280 24 1282 26
rect 1303 43 1305 45
rect 1315 24 1317 26
rect 1337 31 1339 33
rect 1385 31 1387 33
rect 1395 38 1397 40
rect 1395 31 1397 33
rect 1405 33 1407 35
rect 1356 24 1358 26
rect 1448 43 1450 45
rect 1436 24 1438 26
rect 1471 31 1473 33
rect 1471 24 1473 26
rect 1483 39 1485 41
rect 1483 32 1485 34
rect 1493 31 1495 33
rect 1493 24 1495 26
rect 1525 31 1527 33
rect 1525 24 1527 26
rect 1535 39 1537 41
rect 1535 32 1537 34
rect 1547 31 1549 33
rect 1547 24 1549 26
rect 1570 43 1572 45
rect 1582 24 1584 26
rect 1604 31 1606 33
rect 1652 31 1654 33
rect 1662 38 1664 40
rect 1662 31 1664 33
rect 1672 33 1674 35
rect 1623 24 1625 26
rect 1715 43 1717 45
rect 1703 24 1705 26
rect 1738 31 1740 33
rect 1738 24 1740 26
rect 1750 39 1752 41
rect 1750 32 1752 34
rect 1760 31 1762 33
rect 1760 24 1762 26
rect 1792 31 1794 33
rect 1792 24 1794 26
rect 1802 39 1804 41
rect 1802 32 1804 34
rect 1814 31 1816 33
rect 1814 24 1816 26
rect 1837 43 1839 45
rect 1849 24 1851 26
rect 1871 31 1873 33
rect 1922 45 1924 47
rect 1890 24 1892 26
rect 1932 31 1934 33
rect 1948 45 1950 47
rect 1948 38 1950 40
rect 1932 24 1934 26
rect 1968 30 1970 32
rect 2001 43 2003 45
rect 1989 24 1991 26
rect 2024 31 2026 33
rect 2024 24 2026 26
rect 2036 39 2038 41
rect 2036 32 2038 34
rect 2046 31 2048 33
rect 2046 24 2048 26
rect 2078 31 2080 33
rect 2078 24 2080 26
rect 2088 39 2090 41
rect 2088 32 2090 34
rect 2100 31 2102 33
rect 2100 24 2102 26
rect 2123 43 2125 45
rect 2135 24 2137 26
rect 2157 31 2159 33
rect 2201 46 2203 48
rect 2269 46 2271 48
rect 2176 24 2178 26
rect 2211 24 2213 26
rect 2228 34 2230 36
rect 2245 24 2247 26
rect 2279 24 2281 26
rect 2296 34 2298 36
rect 2313 24 2315 26
rect 10 -1 12 1
rect 20 -1 22 1
rect 20 -8 22 -6
rect 30 -3 32 -1
rect 50 -1 52 1
rect 60 -1 62 1
rect 60 -8 62 -6
rect 70 -3 72 -1
rect 101 6 103 8
rect 113 -13 115 -11
rect 136 6 138 8
rect 136 -1 138 1
rect 148 -2 150 0
rect 148 -9 150 -7
rect 158 6 160 8
rect 158 -1 160 1
rect 190 6 192 8
rect 190 -1 192 1
rect 200 -2 202 0
rect 200 -9 202 -7
rect 212 6 214 8
rect 212 -1 214 1
rect 247 6 249 8
rect 235 -13 237 -11
rect 269 -1 271 1
rect 288 6 290 8
rect 317 -1 319 1
rect 327 -1 329 1
rect 327 -8 329 -6
rect 337 -3 339 -1
rect 368 6 370 8
rect 380 -13 382 -11
rect 403 6 405 8
rect 403 -1 405 1
rect 415 -2 417 0
rect 415 -9 417 -7
rect 425 6 427 8
rect 425 -1 427 1
rect 457 6 459 8
rect 457 -1 459 1
rect 467 -2 469 0
rect 467 -9 469 -7
rect 479 6 481 8
rect 479 -1 481 1
rect 514 6 516 8
rect 502 -13 504 -11
rect 536 -1 538 1
rect 555 6 557 8
rect 584 -1 586 1
rect 594 -1 596 1
rect 594 -8 596 -6
rect 604 -3 606 -1
rect 635 6 637 8
rect 647 -13 649 -11
rect 670 6 672 8
rect 670 -1 672 1
rect 682 -2 684 0
rect 682 -9 684 -7
rect 692 6 694 8
rect 692 -1 694 1
rect 724 6 726 8
rect 724 -1 726 1
rect 734 -2 736 0
rect 734 -9 736 -7
rect 746 6 748 8
rect 746 -1 748 1
rect 781 6 783 8
rect 769 -13 771 -11
rect 803 -1 805 1
rect 822 6 824 8
rect 851 -1 853 1
rect 861 -1 863 1
rect 861 -8 863 -6
rect 871 -3 873 -1
rect 902 6 904 8
rect 914 -13 916 -11
rect 937 6 939 8
rect 937 -1 939 1
rect 949 -2 951 0
rect 949 -9 951 -7
rect 959 6 961 8
rect 959 -1 961 1
rect 991 6 993 8
rect 991 -1 993 1
rect 1001 -2 1003 0
rect 1001 -9 1003 -7
rect 1013 6 1015 8
rect 1013 -1 1015 1
rect 1048 6 1050 8
rect 1036 -13 1038 -11
rect 1070 -1 1072 1
rect 1089 6 1091 8
rect 1118 -1 1120 1
rect 1128 -1 1130 1
rect 1128 -8 1130 -6
rect 1138 -3 1140 -1
rect 1169 6 1171 8
rect 1181 -13 1183 -11
rect 1204 6 1206 8
rect 1204 -1 1206 1
rect 1216 -2 1218 0
rect 1216 -9 1218 -7
rect 1226 6 1228 8
rect 1226 -1 1228 1
rect 1258 6 1260 8
rect 1258 -1 1260 1
rect 1268 -2 1270 0
rect 1268 -9 1270 -7
rect 1280 6 1282 8
rect 1280 -1 1282 1
rect 1315 6 1317 8
rect 1303 -13 1305 -11
rect 1337 -1 1339 1
rect 1356 6 1358 8
rect 1385 -1 1387 1
rect 1395 -1 1397 1
rect 1395 -8 1397 -6
rect 1405 -3 1407 -1
rect 1436 6 1438 8
rect 1448 -13 1450 -11
rect 1471 6 1473 8
rect 1471 -1 1473 1
rect 1483 -2 1485 0
rect 1483 -9 1485 -7
rect 1493 6 1495 8
rect 1493 -1 1495 1
rect 1525 6 1527 8
rect 1525 -1 1527 1
rect 1535 -2 1537 0
rect 1535 -9 1537 -7
rect 1547 6 1549 8
rect 1547 -1 1549 1
rect 1582 6 1584 8
rect 1570 -13 1572 -11
rect 1604 -1 1606 1
rect 1623 6 1625 8
rect 1652 -1 1654 1
rect 1662 -1 1664 1
rect 1662 -8 1664 -6
rect 1672 -3 1674 -1
rect 1703 6 1705 8
rect 1715 -13 1717 -11
rect 1738 6 1740 8
rect 1738 -1 1740 1
rect 1750 -2 1752 0
rect 1750 -9 1752 -7
rect 1760 6 1762 8
rect 1760 -1 1762 1
rect 1792 6 1794 8
rect 1792 -1 1794 1
rect 1802 -2 1804 0
rect 1802 -9 1804 -7
rect 1814 6 1816 8
rect 1814 -1 1816 1
rect 1849 6 1851 8
rect 1837 -13 1839 -11
rect 1871 -1 1873 1
rect 1890 6 1892 8
rect 1922 -15 1924 -13
rect 1932 6 1934 8
rect 1932 -1 1934 1
rect 1948 -8 1950 -6
rect 1948 -15 1950 -13
rect 1968 0 1970 2
rect 1989 6 1991 8
rect 2001 -13 2003 -11
rect 2024 6 2026 8
rect 2024 -1 2026 1
rect 2036 -2 2038 0
rect 2036 -9 2038 -7
rect 2046 6 2048 8
rect 2046 -1 2048 1
rect 2078 6 2080 8
rect 2078 -1 2080 1
rect 2088 -2 2090 0
rect 2088 -9 2090 -7
rect 2100 6 2102 8
rect 2100 -1 2102 1
rect 2135 6 2137 8
rect 2123 -13 2125 -11
rect 2157 -1 2159 1
rect 2176 6 2178 8
rect 2211 6 2213 8
rect 2228 -4 2230 -2
rect 2245 6 2247 8
rect 2201 -16 2203 -14
rect 2279 6 2281 8
rect 2296 -4 2298 -2
rect 2313 6 2315 8
rect 2269 -16 2271 -14
rect 10 -113 12 -111
rect 20 -106 22 -104
rect 20 -113 22 -111
rect 30 -111 32 -109
rect 50 -113 52 -111
rect 60 -106 62 -104
rect 60 -113 62 -111
rect 70 -111 72 -109
rect 113 -101 115 -99
rect 101 -120 103 -118
rect 136 -113 138 -111
rect 136 -120 138 -118
rect 148 -105 150 -103
rect 148 -112 150 -110
rect 158 -113 160 -111
rect 158 -120 160 -118
rect 190 -113 192 -111
rect 190 -120 192 -118
rect 200 -105 202 -103
rect 200 -112 202 -110
rect 212 -113 214 -111
rect 212 -120 214 -118
rect 235 -101 237 -99
rect 247 -120 249 -118
rect 269 -113 271 -111
rect 317 -113 319 -111
rect 327 -106 329 -104
rect 327 -113 329 -111
rect 337 -111 339 -109
rect 288 -120 290 -118
rect 380 -101 382 -99
rect 368 -120 370 -118
rect 403 -113 405 -111
rect 403 -120 405 -118
rect 415 -105 417 -103
rect 415 -112 417 -110
rect 425 -113 427 -111
rect 425 -120 427 -118
rect 457 -113 459 -111
rect 457 -120 459 -118
rect 467 -105 469 -103
rect 467 -112 469 -110
rect 479 -113 481 -111
rect 479 -120 481 -118
rect 502 -101 504 -99
rect 514 -120 516 -118
rect 536 -113 538 -111
rect 584 -113 586 -111
rect 594 -106 596 -104
rect 594 -113 596 -111
rect 604 -111 606 -109
rect 555 -120 557 -118
rect 647 -101 649 -99
rect 635 -120 637 -118
rect 670 -113 672 -111
rect 670 -120 672 -118
rect 682 -105 684 -103
rect 682 -112 684 -110
rect 692 -113 694 -111
rect 692 -120 694 -118
rect 724 -113 726 -111
rect 724 -120 726 -118
rect 734 -105 736 -103
rect 734 -112 736 -110
rect 746 -113 748 -111
rect 746 -120 748 -118
rect 769 -101 771 -99
rect 781 -120 783 -118
rect 803 -113 805 -111
rect 851 -113 853 -111
rect 861 -106 863 -104
rect 861 -113 863 -111
rect 871 -111 873 -109
rect 822 -120 824 -118
rect 914 -101 916 -99
rect 902 -120 904 -118
rect 937 -113 939 -111
rect 937 -120 939 -118
rect 949 -105 951 -103
rect 949 -112 951 -110
rect 959 -113 961 -111
rect 959 -120 961 -118
rect 991 -113 993 -111
rect 991 -120 993 -118
rect 1001 -105 1003 -103
rect 1001 -112 1003 -110
rect 1013 -113 1015 -111
rect 1013 -120 1015 -118
rect 1036 -101 1038 -99
rect 1048 -120 1050 -118
rect 1070 -113 1072 -111
rect 1118 -113 1120 -111
rect 1128 -106 1130 -104
rect 1128 -113 1130 -111
rect 1138 -111 1140 -109
rect 1089 -120 1091 -118
rect 1181 -101 1183 -99
rect 1169 -120 1171 -118
rect 1204 -113 1206 -111
rect 1204 -120 1206 -118
rect 1216 -105 1218 -103
rect 1216 -112 1218 -110
rect 1226 -113 1228 -111
rect 1226 -120 1228 -118
rect 1258 -113 1260 -111
rect 1258 -120 1260 -118
rect 1268 -105 1270 -103
rect 1268 -112 1270 -110
rect 1280 -113 1282 -111
rect 1280 -120 1282 -118
rect 1303 -101 1305 -99
rect 1315 -120 1317 -118
rect 1337 -113 1339 -111
rect 1385 -113 1387 -111
rect 1395 -106 1397 -104
rect 1395 -113 1397 -111
rect 1405 -111 1407 -109
rect 1356 -120 1358 -118
rect 1448 -101 1450 -99
rect 1436 -120 1438 -118
rect 1471 -113 1473 -111
rect 1471 -120 1473 -118
rect 1483 -105 1485 -103
rect 1483 -112 1485 -110
rect 1493 -113 1495 -111
rect 1493 -120 1495 -118
rect 1525 -113 1527 -111
rect 1525 -120 1527 -118
rect 1535 -105 1537 -103
rect 1535 -112 1537 -110
rect 1547 -113 1549 -111
rect 1547 -120 1549 -118
rect 1570 -101 1572 -99
rect 1582 -120 1584 -118
rect 1604 -113 1606 -111
rect 1652 -113 1654 -111
rect 1662 -106 1664 -104
rect 1662 -113 1664 -111
rect 1672 -111 1674 -109
rect 1623 -120 1625 -118
rect 1715 -101 1717 -99
rect 1703 -120 1705 -118
rect 1738 -113 1740 -111
rect 1738 -120 1740 -118
rect 1750 -105 1752 -103
rect 1750 -112 1752 -110
rect 1760 -113 1762 -111
rect 1760 -120 1762 -118
rect 1792 -113 1794 -111
rect 1792 -120 1794 -118
rect 1802 -105 1804 -103
rect 1802 -112 1804 -110
rect 1814 -113 1816 -111
rect 1814 -120 1816 -118
rect 1837 -101 1839 -99
rect 1849 -120 1851 -118
rect 1871 -113 1873 -111
rect 1922 -99 1924 -97
rect 1890 -120 1892 -118
rect 1932 -113 1934 -111
rect 1948 -99 1950 -97
rect 1948 -106 1950 -104
rect 1932 -120 1934 -118
rect 1968 -114 1970 -112
rect 2001 -101 2003 -99
rect 1989 -120 1991 -118
rect 2024 -113 2026 -111
rect 2024 -120 2026 -118
rect 2036 -105 2038 -103
rect 2036 -112 2038 -110
rect 2046 -113 2048 -111
rect 2046 -120 2048 -118
rect 2078 -113 2080 -111
rect 2078 -120 2080 -118
rect 2088 -105 2090 -103
rect 2088 -112 2090 -110
rect 2100 -113 2102 -111
rect 2100 -120 2102 -118
rect 2123 -101 2125 -99
rect 2135 -120 2137 -118
rect 2157 -113 2159 -111
rect 2201 -98 2203 -96
rect 2269 -98 2271 -96
rect 2176 -120 2178 -118
rect 2211 -120 2213 -118
rect 2228 -110 2230 -108
rect 2245 -120 2247 -118
rect 2279 -120 2281 -118
rect 2296 -110 2298 -108
rect 2313 -120 2315 -118
rect 10 -145 12 -143
rect 20 -145 22 -143
rect 20 -152 22 -150
rect 30 -147 32 -145
rect 50 -145 52 -143
rect 60 -145 62 -143
rect 60 -152 62 -150
rect 70 -147 72 -145
rect 101 -138 103 -136
rect 113 -157 115 -155
rect 136 -138 138 -136
rect 136 -145 138 -143
rect 148 -146 150 -144
rect 148 -153 150 -151
rect 158 -138 160 -136
rect 158 -145 160 -143
rect 190 -138 192 -136
rect 190 -145 192 -143
rect 200 -146 202 -144
rect 200 -153 202 -151
rect 212 -138 214 -136
rect 212 -145 214 -143
rect 247 -138 249 -136
rect 235 -157 237 -155
rect 269 -145 271 -143
rect 288 -138 290 -136
rect 317 -145 319 -143
rect 327 -145 329 -143
rect 327 -152 329 -150
rect 337 -147 339 -145
rect 368 -138 370 -136
rect 380 -157 382 -155
rect 403 -138 405 -136
rect 403 -145 405 -143
rect 415 -146 417 -144
rect 415 -153 417 -151
rect 425 -138 427 -136
rect 425 -145 427 -143
rect 457 -138 459 -136
rect 457 -145 459 -143
rect 467 -146 469 -144
rect 467 -153 469 -151
rect 479 -138 481 -136
rect 479 -145 481 -143
rect 514 -138 516 -136
rect 502 -157 504 -155
rect 536 -145 538 -143
rect 555 -138 557 -136
rect 584 -145 586 -143
rect 594 -145 596 -143
rect 594 -152 596 -150
rect 604 -147 606 -145
rect 635 -138 637 -136
rect 647 -157 649 -155
rect 670 -138 672 -136
rect 670 -145 672 -143
rect 682 -146 684 -144
rect 682 -153 684 -151
rect 692 -138 694 -136
rect 692 -145 694 -143
rect 724 -138 726 -136
rect 724 -145 726 -143
rect 734 -146 736 -144
rect 734 -153 736 -151
rect 746 -138 748 -136
rect 746 -145 748 -143
rect 781 -138 783 -136
rect 769 -157 771 -155
rect 803 -145 805 -143
rect 822 -138 824 -136
rect 851 -145 853 -143
rect 861 -145 863 -143
rect 861 -152 863 -150
rect 871 -147 873 -145
rect 902 -138 904 -136
rect 914 -157 916 -155
rect 937 -138 939 -136
rect 937 -145 939 -143
rect 949 -146 951 -144
rect 949 -153 951 -151
rect 959 -138 961 -136
rect 959 -145 961 -143
rect 991 -138 993 -136
rect 991 -145 993 -143
rect 1001 -146 1003 -144
rect 1001 -153 1003 -151
rect 1013 -138 1015 -136
rect 1013 -145 1015 -143
rect 1048 -138 1050 -136
rect 1036 -157 1038 -155
rect 1070 -145 1072 -143
rect 1089 -138 1091 -136
rect 1118 -145 1120 -143
rect 1128 -145 1130 -143
rect 1128 -152 1130 -150
rect 1138 -147 1140 -145
rect 1169 -138 1171 -136
rect 1181 -157 1183 -155
rect 1204 -138 1206 -136
rect 1204 -145 1206 -143
rect 1216 -146 1218 -144
rect 1216 -153 1218 -151
rect 1226 -138 1228 -136
rect 1226 -145 1228 -143
rect 1258 -138 1260 -136
rect 1258 -145 1260 -143
rect 1268 -146 1270 -144
rect 1268 -153 1270 -151
rect 1280 -138 1282 -136
rect 1280 -145 1282 -143
rect 1315 -138 1317 -136
rect 1303 -157 1305 -155
rect 1337 -145 1339 -143
rect 1356 -138 1358 -136
rect 1385 -145 1387 -143
rect 1395 -145 1397 -143
rect 1395 -152 1397 -150
rect 1405 -147 1407 -145
rect 1436 -138 1438 -136
rect 1448 -157 1450 -155
rect 1471 -138 1473 -136
rect 1471 -145 1473 -143
rect 1483 -146 1485 -144
rect 1483 -153 1485 -151
rect 1493 -138 1495 -136
rect 1493 -145 1495 -143
rect 1525 -138 1527 -136
rect 1525 -145 1527 -143
rect 1535 -146 1537 -144
rect 1535 -153 1537 -151
rect 1547 -138 1549 -136
rect 1547 -145 1549 -143
rect 1582 -138 1584 -136
rect 1570 -157 1572 -155
rect 1604 -145 1606 -143
rect 1623 -138 1625 -136
rect 1652 -145 1654 -143
rect 1662 -145 1664 -143
rect 1662 -152 1664 -150
rect 1672 -147 1674 -145
rect 1703 -138 1705 -136
rect 1715 -157 1717 -155
rect 1738 -138 1740 -136
rect 1738 -145 1740 -143
rect 1750 -146 1752 -144
rect 1750 -153 1752 -151
rect 1760 -138 1762 -136
rect 1760 -145 1762 -143
rect 1792 -138 1794 -136
rect 1792 -145 1794 -143
rect 1802 -146 1804 -144
rect 1802 -153 1804 -151
rect 1814 -138 1816 -136
rect 1814 -145 1816 -143
rect 1849 -138 1851 -136
rect 1837 -157 1839 -155
rect 1871 -145 1873 -143
rect 1890 -138 1892 -136
rect 1922 -159 1924 -157
rect 1932 -138 1934 -136
rect 1932 -145 1934 -143
rect 1948 -152 1950 -150
rect 1948 -159 1950 -157
rect 1968 -144 1970 -142
rect 1989 -138 1991 -136
rect 2001 -157 2003 -155
rect 2024 -138 2026 -136
rect 2024 -145 2026 -143
rect 2036 -146 2038 -144
rect 2036 -153 2038 -151
rect 2046 -138 2048 -136
rect 2046 -145 2048 -143
rect 2078 -138 2080 -136
rect 2078 -145 2080 -143
rect 2088 -146 2090 -144
rect 2088 -153 2090 -151
rect 2100 -138 2102 -136
rect 2100 -145 2102 -143
rect 2135 -138 2137 -136
rect 2123 -157 2125 -155
rect 2157 -145 2159 -143
rect 2176 -138 2178 -136
rect 2211 -138 2213 -136
rect 2228 -148 2230 -146
rect 2245 -138 2247 -136
rect 2201 -160 2203 -158
rect 2279 -138 2281 -136
rect 2296 -148 2298 -146
rect 2313 -138 2315 -136
rect 2269 -160 2271 -158
rect 10 -257 12 -255
rect 20 -250 22 -248
rect 20 -257 22 -255
rect 30 -255 32 -253
rect 50 -257 52 -255
rect 60 -250 62 -248
rect 60 -257 62 -255
rect 70 -255 72 -253
rect 113 -245 115 -243
rect 101 -264 103 -262
rect 136 -257 138 -255
rect 136 -264 138 -262
rect 148 -249 150 -247
rect 148 -256 150 -254
rect 158 -257 160 -255
rect 158 -264 160 -262
rect 190 -257 192 -255
rect 190 -264 192 -262
rect 200 -249 202 -247
rect 200 -256 202 -254
rect 212 -257 214 -255
rect 212 -264 214 -262
rect 235 -245 237 -243
rect 247 -264 249 -262
rect 269 -257 271 -255
rect 317 -257 319 -255
rect 327 -250 329 -248
rect 327 -257 329 -255
rect 337 -255 339 -253
rect 288 -264 290 -262
rect 380 -245 382 -243
rect 368 -264 370 -262
rect 403 -257 405 -255
rect 403 -264 405 -262
rect 415 -249 417 -247
rect 415 -256 417 -254
rect 425 -257 427 -255
rect 425 -264 427 -262
rect 457 -257 459 -255
rect 457 -264 459 -262
rect 467 -249 469 -247
rect 467 -256 469 -254
rect 479 -257 481 -255
rect 479 -264 481 -262
rect 502 -245 504 -243
rect 514 -264 516 -262
rect 536 -257 538 -255
rect 584 -257 586 -255
rect 594 -250 596 -248
rect 594 -257 596 -255
rect 604 -255 606 -253
rect 555 -264 557 -262
rect 647 -245 649 -243
rect 635 -264 637 -262
rect 670 -257 672 -255
rect 670 -264 672 -262
rect 682 -249 684 -247
rect 682 -256 684 -254
rect 692 -257 694 -255
rect 692 -264 694 -262
rect 724 -257 726 -255
rect 724 -264 726 -262
rect 734 -249 736 -247
rect 734 -256 736 -254
rect 746 -257 748 -255
rect 746 -264 748 -262
rect 769 -245 771 -243
rect 781 -264 783 -262
rect 803 -257 805 -255
rect 851 -257 853 -255
rect 861 -250 863 -248
rect 861 -257 863 -255
rect 871 -255 873 -253
rect 822 -264 824 -262
rect 914 -245 916 -243
rect 902 -264 904 -262
rect 937 -257 939 -255
rect 937 -264 939 -262
rect 949 -249 951 -247
rect 949 -256 951 -254
rect 959 -257 961 -255
rect 959 -264 961 -262
rect 991 -257 993 -255
rect 991 -264 993 -262
rect 1001 -249 1003 -247
rect 1001 -256 1003 -254
rect 1013 -257 1015 -255
rect 1013 -264 1015 -262
rect 1036 -245 1038 -243
rect 1048 -264 1050 -262
rect 1070 -257 1072 -255
rect 1118 -257 1120 -255
rect 1128 -250 1130 -248
rect 1128 -257 1130 -255
rect 1138 -255 1140 -253
rect 1089 -264 1091 -262
rect 1181 -245 1183 -243
rect 1169 -264 1171 -262
rect 1204 -257 1206 -255
rect 1204 -264 1206 -262
rect 1216 -249 1218 -247
rect 1216 -256 1218 -254
rect 1226 -257 1228 -255
rect 1226 -264 1228 -262
rect 1258 -257 1260 -255
rect 1258 -264 1260 -262
rect 1268 -249 1270 -247
rect 1268 -256 1270 -254
rect 1280 -257 1282 -255
rect 1280 -264 1282 -262
rect 1303 -245 1305 -243
rect 1315 -264 1317 -262
rect 1337 -257 1339 -255
rect 1385 -257 1387 -255
rect 1395 -250 1397 -248
rect 1395 -257 1397 -255
rect 1405 -255 1407 -253
rect 1356 -264 1358 -262
rect 1448 -245 1450 -243
rect 1436 -264 1438 -262
rect 1471 -257 1473 -255
rect 1471 -264 1473 -262
rect 1483 -249 1485 -247
rect 1483 -256 1485 -254
rect 1493 -257 1495 -255
rect 1493 -264 1495 -262
rect 1525 -257 1527 -255
rect 1525 -264 1527 -262
rect 1535 -249 1537 -247
rect 1535 -256 1537 -254
rect 1547 -257 1549 -255
rect 1547 -264 1549 -262
rect 1570 -245 1572 -243
rect 1582 -264 1584 -262
rect 1604 -257 1606 -255
rect 1652 -257 1654 -255
rect 1662 -250 1664 -248
rect 1662 -257 1664 -255
rect 1672 -255 1674 -253
rect 1623 -264 1625 -262
rect 1715 -245 1717 -243
rect 1703 -264 1705 -262
rect 1738 -257 1740 -255
rect 1738 -264 1740 -262
rect 1750 -249 1752 -247
rect 1750 -256 1752 -254
rect 1760 -257 1762 -255
rect 1760 -264 1762 -262
rect 1792 -257 1794 -255
rect 1792 -264 1794 -262
rect 1802 -249 1804 -247
rect 1802 -256 1804 -254
rect 1814 -257 1816 -255
rect 1814 -264 1816 -262
rect 1837 -245 1839 -243
rect 1849 -264 1851 -262
rect 1871 -257 1873 -255
rect 1922 -243 1924 -241
rect 1890 -264 1892 -262
rect 1932 -257 1934 -255
rect 1948 -243 1950 -241
rect 1948 -250 1950 -248
rect 1932 -264 1934 -262
rect 1968 -258 1970 -256
rect 2001 -245 2003 -243
rect 1989 -264 1991 -262
rect 2024 -257 2026 -255
rect 2024 -264 2026 -262
rect 2036 -249 2038 -247
rect 2036 -256 2038 -254
rect 2046 -257 2048 -255
rect 2046 -264 2048 -262
rect 2078 -257 2080 -255
rect 2078 -264 2080 -262
rect 2088 -249 2090 -247
rect 2088 -256 2090 -254
rect 2100 -257 2102 -255
rect 2100 -264 2102 -262
rect 2123 -245 2125 -243
rect 2135 -264 2137 -262
rect 2157 -257 2159 -255
rect 2201 -242 2203 -240
rect 2269 -242 2271 -240
rect 2176 -264 2178 -262
rect 2211 -264 2213 -262
rect 2228 -254 2230 -252
rect 2245 -264 2247 -262
rect 2279 -264 2281 -262
rect 2296 -254 2298 -252
rect 2313 -264 2315 -262
<< pdifct1 >>
rect 40 280 42 282
rect 40 273 42 275
rect 80 280 82 282
rect 80 273 82 275
rect 90 282 92 284
rect 90 275 92 277
rect 168 279 170 281
rect 168 272 170 274
rect 180 279 182 281
rect 180 272 182 274
rect 258 282 260 284
rect 258 275 260 277
rect 299 284 301 286
rect 299 277 301 279
rect 347 280 349 282
rect 347 273 349 275
rect 357 282 359 284
rect 357 275 359 277
rect 435 279 437 281
rect 435 272 437 274
rect 447 279 449 281
rect 447 272 449 274
rect 525 282 527 284
rect 525 275 527 277
rect 566 284 568 286
rect 566 277 568 279
rect 614 280 616 282
rect 614 273 616 275
rect 624 282 626 284
rect 624 275 626 277
rect 702 279 704 281
rect 702 272 704 274
rect 714 279 716 281
rect 714 272 716 274
rect 792 282 794 284
rect 792 275 794 277
rect 833 284 835 286
rect 833 277 835 279
rect 881 280 883 282
rect 881 273 883 275
rect 891 282 893 284
rect 891 275 893 277
rect 969 279 971 281
rect 969 272 971 274
rect 981 279 983 281
rect 981 272 983 274
rect 1059 282 1061 284
rect 1059 275 1061 277
rect 1100 284 1102 286
rect 1100 277 1102 279
rect 1148 280 1150 282
rect 1148 273 1150 275
rect 1158 282 1160 284
rect 1158 275 1160 277
rect 1236 279 1238 281
rect 1236 272 1238 274
rect 1248 279 1250 281
rect 1248 272 1250 274
rect 1326 282 1328 284
rect 1326 275 1328 277
rect 1367 284 1369 286
rect 1367 277 1369 279
rect 1415 280 1417 282
rect 1415 273 1417 275
rect 1425 282 1427 284
rect 1425 275 1427 277
rect 1503 279 1505 281
rect 1503 272 1505 274
rect 1515 279 1517 281
rect 1515 272 1517 274
rect 1593 282 1595 284
rect 1593 275 1595 277
rect 1634 284 1636 286
rect 1634 277 1636 279
rect 1682 280 1684 282
rect 1682 273 1684 275
rect 1692 282 1694 284
rect 1692 275 1694 277
rect 1770 279 1772 281
rect 1770 272 1772 274
rect 1782 279 1784 281
rect 1782 272 1784 274
rect 1860 282 1862 284
rect 1860 275 1862 277
rect 1901 284 1903 286
rect 1901 277 1903 279
rect 1958 280 1960 282
rect 1978 282 1980 284
rect 1978 275 1980 277
rect 2056 279 2058 281
rect 2056 272 2058 274
rect 2068 279 2070 281
rect 2068 272 2070 274
rect 2146 282 2148 284
rect 2146 275 2148 277
rect 2187 284 2189 286
rect 2187 277 2189 279
rect 2255 287 2257 289
rect 2323 287 2325 289
rect 40 188 42 190
rect 40 180 42 182
rect 80 189 82 191
rect 80 182 82 184
rect 90 187 92 189
rect 90 180 92 182
rect 168 190 170 192
rect 168 183 170 185
rect 180 190 182 192
rect 180 183 182 185
rect 258 187 260 189
rect 258 180 260 182
rect 299 185 301 187
rect 299 178 301 180
rect 347 189 349 191
rect 347 182 349 184
rect 357 187 359 189
rect 357 180 359 182
rect 435 190 437 192
rect 435 183 437 185
rect 447 190 449 192
rect 447 183 449 185
rect 525 187 527 189
rect 525 180 527 182
rect 566 185 568 187
rect 566 178 568 180
rect 614 189 616 191
rect 614 182 616 184
rect 624 187 626 189
rect 624 180 626 182
rect 702 190 704 192
rect 702 183 704 185
rect 714 190 716 192
rect 714 183 716 185
rect 792 187 794 189
rect 792 180 794 182
rect 833 185 835 187
rect 833 178 835 180
rect 881 189 883 191
rect 881 182 883 184
rect 891 187 893 189
rect 891 180 893 182
rect 969 190 971 192
rect 969 183 971 185
rect 981 190 983 192
rect 981 183 983 185
rect 1059 187 1061 189
rect 1059 180 1061 182
rect 1100 185 1102 187
rect 1100 178 1102 180
rect 1148 189 1150 191
rect 1148 182 1150 184
rect 1158 187 1160 189
rect 1158 180 1160 182
rect 1236 190 1238 192
rect 1236 183 1238 185
rect 1248 190 1250 192
rect 1248 183 1250 185
rect 1326 187 1328 189
rect 1326 180 1328 182
rect 1367 185 1369 187
rect 1367 178 1369 180
rect 1415 189 1417 191
rect 1415 182 1417 184
rect 1425 187 1427 189
rect 1425 180 1427 182
rect 1503 190 1505 192
rect 1503 183 1505 185
rect 1515 190 1517 192
rect 1515 183 1517 185
rect 1593 187 1595 189
rect 1593 180 1595 182
rect 1634 185 1636 187
rect 1634 178 1636 180
rect 1682 189 1684 191
rect 1682 182 1684 184
rect 1692 187 1694 189
rect 1692 180 1694 182
rect 1770 190 1772 192
rect 1770 183 1772 185
rect 1782 190 1784 192
rect 1782 183 1784 185
rect 1860 187 1862 189
rect 1860 180 1862 182
rect 1901 185 1903 187
rect 1901 178 1903 180
rect 1958 182 1960 184
rect 1978 187 1980 189
rect 1978 180 1980 182
rect 2056 190 2058 192
rect 2056 183 2058 185
rect 2068 190 2070 192
rect 2068 183 2070 185
rect 2146 187 2148 189
rect 2146 180 2148 182
rect 2187 185 2189 187
rect 2187 178 2189 180
rect 2255 175 2257 177
rect 2323 175 2325 177
rect 40 139 42 141
rect 40 131 42 133
rect 80 136 82 138
rect 80 129 82 131
rect 90 138 92 140
rect 90 131 92 133
rect 168 135 170 137
rect 168 128 170 130
rect 180 135 182 137
rect 180 128 182 130
rect 258 138 260 140
rect 258 131 260 133
rect 299 140 301 142
rect 299 133 301 135
rect 347 136 349 138
rect 347 129 349 131
rect 357 138 359 140
rect 357 131 359 133
rect 435 135 437 137
rect 435 128 437 130
rect 447 135 449 137
rect 447 128 449 130
rect 525 138 527 140
rect 525 131 527 133
rect 566 140 568 142
rect 566 133 568 135
rect 614 136 616 138
rect 614 129 616 131
rect 624 138 626 140
rect 624 131 626 133
rect 702 135 704 137
rect 702 128 704 130
rect 714 135 716 137
rect 714 128 716 130
rect 792 138 794 140
rect 792 131 794 133
rect 833 140 835 142
rect 833 133 835 135
rect 881 136 883 138
rect 881 129 883 131
rect 891 138 893 140
rect 891 131 893 133
rect 969 135 971 137
rect 969 128 971 130
rect 981 135 983 137
rect 981 128 983 130
rect 1059 138 1061 140
rect 1059 131 1061 133
rect 1100 140 1102 142
rect 1100 133 1102 135
rect 1148 136 1150 138
rect 1148 129 1150 131
rect 1158 138 1160 140
rect 1158 131 1160 133
rect 1236 135 1238 137
rect 1236 128 1238 130
rect 1248 135 1250 137
rect 1248 128 1250 130
rect 1326 138 1328 140
rect 1326 131 1328 133
rect 1367 140 1369 142
rect 1367 133 1369 135
rect 1415 136 1417 138
rect 1415 129 1417 131
rect 1425 138 1427 140
rect 1425 131 1427 133
rect 1503 135 1505 137
rect 1503 128 1505 130
rect 1515 135 1517 137
rect 1515 128 1517 130
rect 1593 138 1595 140
rect 1593 131 1595 133
rect 1634 140 1636 142
rect 1634 133 1636 135
rect 1682 136 1684 138
rect 1682 129 1684 131
rect 1692 138 1694 140
rect 1692 131 1694 133
rect 1770 135 1772 137
rect 1770 128 1772 130
rect 1782 135 1784 137
rect 1782 128 1784 130
rect 1860 138 1862 140
rect 1860 131 1862 133
rect 1901 140 1903 142
rect 1901 133 1903 135
rect 1958 136 1960 138
rect 1978 138 1980 140
rect 1978 131 1980 133
rect 2056 135 2058 137
rect 2056 128 2058 130
rect 2068 135 2070 137
rect 2068 128 2070 130
rect 2146 138 2148 140
rect 2146 131 2148 133
rect 2187 140 2189 142
rect 2187 133 2189 135
rect 2255 143 2257 145
rect 2323 143 2325 145
rect 40 42 42 44
rect 40 35 42 37
rect 80 45 82 47
rect 80 38 82 40
rect 90 43 92 45
rect 90 36 92 38
rect 168 46 170 48
rect 168 39 170 41
rect 180 46 182 48
rect 180 39 182 41
rect 258 43 260 45
rect 258 36 260 38
rect 299 41 301 43
rect 299 34 301 36
rect 347 45 349 47
rect 347 38 349 40
rect 357 43 359 45
rect 357 36 359 38
rect 435 46 437 48
rect 435 39 437 41
rect 447 46 449 48
rect 447 39 449 41
rect 525 43 527 45
rect 525 36 527 38
rect 566 41 568 43
rect 566 34 568 36
rect 614 45 616 47
rect 614 38 616 40
rect 624 43 626 45
rect 624 36 626 38
rect 702 46 704 48
rect 702 39 704 41
rect 714 46 716 48
rect 714 39 716 41
rect 792 43 794 45
rect 792 36 794 38
rect 833 41 835 43
rect 833 34 835 36
rect 881 45 883 47
rect 881 38 883 40
rect 891 43 893 45
rect 891 36 893 38
rect 969 46 971 48
rect 969 39 971 41
rect 981 46 983 48
rect 981 39 983 41
rect 1059 43 1061 45
rect 1059 36 1061 38
rect 1100 41 1102 43
rect 1100 34 1102 36
rect 1148 45 1150 47
rect 1148 38 1150 40
rect 1158 43 1160 45
rect 1158 36 1160 38
rect 1236 46 1238 48
rect 1236 39 1238 41
rect 1248 46 1250 48
rect 1248 39 1250 41
rect 1326 43 1328 45
rect 1326 36 1328 38
rect 1367 41 1369 43
rect 1367 34 1369 36
rect 1415 45 1417 47
rect 1415 38 1417 40
rect 1425 43 1427 45
rect 1425 36 1427 38
rect 1503 46 1505 48
rect 1503 39 1505 41
rect 1515 46 1517 48
rect 1515 39 1517 41
rect 1593 43 1595 45
rect 1593 36 1595 38
rect 1634 41 1636 43
rect 1634 34 1636 36
rect 1682 45 1684 47
rect 1682 38 1684 40
rect 1692 43 1694 45
rect 1692 36 1694 38
rect 1770 46 1772 48
rect 1770 39 1772 41
rect 1782 46 1784 48
rect 1782 39 1784 41
rect 1860 43 1862 45
rect 1860 36 1862 38
rect 1901 41 1903 43
rect 1901 34 1903 36
rect 1958 38 1960 40
rect 1978 43 1980 45
rect 1978 36 1980 38
rect 2056 46 2058 48
rect 2056 39 2058 41
rect 2068 46 2070 48
rect 2068 39 2070 41
rect 2146 43 2148 45
rect 2146 36 2148 38
rect 2187 41 2189 43
rect 2187 34 2189 36
rect 2255 31 2257 33
rect 2323 31 2325 33
rect 40 -8 42 -6
rect 40 -15 42 -13
rect 80 -8 82 -6
rect 80 -15 82 -13
rect 90 -6 92 -4
rect 90 -13 92 -11
rect 168 -9 170 -7
rect 168 -16 170 -14
rect 180 -9 182 -7
rect 180 -16 182 -14
rect 258 -6 260 -4
rect 258 -13 260 -11
rect 299 -4 301 -2
rect 299 -11 301 -9
rect 347 -8 349 -6
rect 347 -15 349 -13
rect 357 -6 359 -4
rect 357 -13 359 -11
rect 435 -9 437 -7
rect 435 -16 437 -14
rect 447 -9 449 -7
rect 447 -16 449 -14
rect 525 -6 527 -4
rect 525 -13 527 -11
rect 566 -4 568 -2
rect 566 -11 568 -9
rect 614 -8 616 -6
rect 614 -15 616 -13
rect 624 -6 626 -4
rect 624 -13 626 -11
rect 702 -9 704 -7
rect 702 -16 704 -14
rect 714 -9 716 -7
rect 714 -16 716 -14
rect 792 -6 794 -4
rect 792 -13 794 -11
rect 833 -4 835 -2
rect 833 -11 835 -9
rect 881 -8 883 -6
rect 881 -15 883 -13
rect 891 -6 893 -4
rect 891 -13 893 -11
rect 969 -9 971 -7
rect 969 -16 971 -14
rect 981 -9 983 -7
rect 981 -16 983 -14
rect 1059 -6 1061 -4
rect 1059 -13 1061 -11
rect 1100 -4 1102 -2
rect 1100 -11 1102 -9
rect 1148 -8 1150 -6
rect 1148 -15 1150 -13
rect 1158 -6 1160 -4
rect 1158 -13 1160 -11
rect 1236 -9 1238 -7
rect 1236 -16 1238 -14
rect 1248 -9 1250 -7
rect 1248 -16 1250 -14
rect 1326 -6 1328 -4
rect 1326 -13 1328 -11
rect 1367 -4 1369 -2
rect 1367 -11 1369 -9
rect 1415 -8 1417 -6
rect 1415 -15 1417 -13
rect 1425 -6 1427 -4
rect 1425 -13 1427 -11
rect 1503 -9 1505 -7
rect 1503 -16 1505 -14
rect 1515 -9 1517 -7
rect 1515 -16 1517 -14
rect 1593 -6 1595 -4
rect 1593 -13 1595 -11
rect 1634 -4 1636 -2
rect 1634 -11 1636 -9
rect 1682 -8 1684 -6
rect 1682 -15 1684 -13
rect 1692 -6 1694 -4
rect 1692 -13 1694 -11
rect 1770 -9 1772 -7
rect 1770 -16 1772 -14
rect 1782 -9 1784 -7
rect 1782 -16 1784 -14
rect 1860 -6 1862 -4
rect 1860 -13 1862 -11
rect 1901 -4 1903 -2
rect 1901 -11 1903 -9
rect 1958 -8 1960 -6
rect 1978 -6 1980 -4
rect 1978 -13 1980 -11
rect 2056 -9 2058 -7
rect 2056 -16 2058 -14
rect 2068 -9 2070 -7
rect 2068 -16 2070 -14
rect 2146 -6 2148 -4
rect 2146 -13 2148 -11
rect 2187 -4 2189 -2
rect 2187 -11 2189 -9
rect 2255 -1 2257 1
rect 2323 -1 2325 1
rect 40 -100 42 -98
rect 40 -108 42 -106
rect 80 -99 82 -97
rect 80 -106 82 -104
rect 90 -101 92 -99
rect 90 -108 92 -106
rect 168 -98 170 -96
rect 168 -105 170 -103
rect 180 -98 182 -96
rect 180 -105 182 -103
rect 258 -101 260 -99
rect 258 -108 260 -106
rect 299 -103 301 -101
rect 299 -110 301 -108
rect 347 -99 349 -97
rect 347 -106 349 -104
rect 357 -101 359 -99
rect 357 -108 359 -106
rect 435 -98 437 -96
rect 435 -105 437 -103
rect 447 -98 449 -96
rect 447 -105 449 -103
rect 525 -101 527 -99
rect 525 -108 527 -106
rect 566 -103 568 -101
rect 566 -110 568 -108
rect 614 -99 616 -97
rect 614 -106 616 -104
rect 624 -101 626 -99
rect 624 -108 626 -106
rect 702 -98 704 -96
rect 702 -105 704 -103
rect 714 -98 716 -96
rect 714 -105 716 -103
rect 792 -101 794 -99
rect 792 -108 794 -106
rect 833 -103 835 -101
rect 833 -110 835 -108
rect 881 -99 883 -97
rect 881 -106 883 -104
rect 891 -101 893 -99
rect 891 -108 893 -106
rect 969 -98 971 -96
rect 969 -105 971 -103
rect 981 -98 983 -96
rect 981 -105 983 -103
rect 1059 -101 1061 -99
rect 1059 -108 1061 -106
rect 1100 -103 1102 -101
rect 1100 -110 1102 -108
rect 1148 -99 1150 -97
rect 1148 -106 1150 -104
rect 1158 -101 1160 -99
rect 1158 -108 1160 -106
rect 1236 -98 1238 -96
rect 1236 -105 1238 -103
rect 1248 -98 1250 -96
rect 1248 -105 1250 -103
rect 1326 -101 1328 -99
rect 1326 -108 1328 -106
rect 1367 -103 1369 -101
rect 1367 -110 1369 -108
rect 1415 -99 1417 -97
rect 1415 -106 1417 -104
rect 1425 -101 1427 -99
rect 1425 -108 1427 -106
rect 1503 -98 1505 -96
rect 1503 -105 1505 -103
rect 1515 -98 1517 -96
rect 1515 -105 1517 -103
rect 1593 -101 1595 -99
rect 1593 -108 1595 -106
rect 1634 -103 1636 -101
rect 1634 -110 1636 -108
rect 1682 -99 1684 -97
rect 1682 -106 1684 -104
rect 1692 -101 1694 -99
rect 1692 -108 1694 -106
rect 1770 -98 1772 -96
rect 1770 -105 1772 -103
rect 1782 -98 1784 -96
rect 1782 -105 1784 -103
rect 1860 -101 1862 -99
rect 1860 -108 1862 -106
rect 1901 -103 1903 -101
rect 1901 -110 1903 -108
rect 1958 -106 1960 -104
rect 1978 -101 1980 -99
rect 1978 -108 1980 -106
rect 2056 -98 2058 -96
rect 2056 -105 2058 -103
rect 2068 -98 2070 -96
rect 2068 -105 2070 -103
rect 2146 -101 2148 -99
rect 2146 -108 2148 -106
rect 2187 -103 2189 -101
rect 2187 -110 2189 -108
rect 2255 -113 2257 -111
rect 2323 -113 2325 -111
rect 40 -149 42 -147
rect 40 -157 42 -155
rect 80 -152 82 -150
rect 80 -159 82 -157
rect 90 -150 92 -148
rect 90 -157 92 -155
rect 168 -153 170 -151
rect 168 -160 170 -158
rect 180 -153 182 -151
rect 180 -160 182 -158
rect 258 -150 260 -148
rect 258 -157 260 -155
rect 299 -148 301 -146
rect 299 -155 301 -153
rect 347 -152 349 -150
rect 347 -159 349 -157
rect 357 -150 359 -148
rect 357 -157 359 -155
rect 435 -153 437 -151
rect 435 -160 437 -158
rect 447 -153 449 -151
rect 447 -160 449 -158
rect 525 -150 527 -148
rect 525 -157 527 -155
rect 566 -148 568 -146
rect 566 -155 568 -153
rect 614 -152 616 -150
rect 614 -159 616 -157
rect 624 -150 626 -148
rect 624 -157 626 -155
rect 702 -153 704 -151
rect 702 -160 704 -158
rect 714 -153 716 -151
rect 714 -160 716 -158
rect 792 -150 794 -148
rect 792 -157 794 -155
rect 833 -148 835 -146
rect 833 -155 835 -153
rect 881 -152 883 -150
rect 881 -159 883 -157
rect 891 -150 893 -148
rect 891 -157 893 -155
rect 969 -153 971 -151
rect 969 -160 971 -158
rect 981 -153 983 -151
rect 981 -160 983 -158
rect 1059 -150 1061 -148
rect 1059 -157 1061 -155
rect 1100 -148 1102 -146
rect 1100 -155 1102 -153
rect 1148 -152 1150 -150
rect 1148 -159 1150 -157
rect 1158 -150 1160 -148
rect 1158 -157 1160 -155
rect 1236 -153 1238 -151
rect 1236 -160 1238 -158
rect 1248 -153 1250 -151
rect 1248 -160 1250 -158
rect 1326 -150 1328 -148
rect 1326 -157 1328 -155
rect 1367 -148 1369 -146
rect 1367 -155 1369 -153
rect 1415 -152 1417 -150
rect 1415 -159 1417 -157
rect 1425 -150 1427 -148
rect 1425 -157 1427 -155
rect 1503 -153 1505 -151
rect 1503 -160 1505 -158
rect 1515 -153 1517 -151
rect 1515 -160 1517 -158
rect 1593 -150 1595 -148
rect 1593 -157 1595 -155
rect 1634 -148 1636 -146
rect 1634 -155 1636 -153
rect 1682 -152 1684 -150
rect 1682 -159 1684 -157
rect 1692 -150 1694 -148
rect 1692 -157 1694 -155
rect 1770 -153 1772 -151
rect 1770 -160 1772 -158
rect 1782 -153 1784 -151
rect 1782 -160 1784 -158
rect 1860 -150 1862 -148
rect 1860 -157 1862 -155
rect 1901 -148 1903 -146
rect 1901 -155 1903 -153
rect 1958 -152 1960 -150
rect 1978 -150 1980 -148
rect 1978 -157 1980 -155
rect 2056 -153 2058 -151
rect 2056 -160 2058 -158
rect 2068 -153 2070 -151
rect 2068 -160 2070 -158
rect 2146 -150 2148 -148
rect 2146 -157 2148 -155
rect 2187 -148 2189 -146
rect 2187 -155 2189 -153
rect 2255 -145 2257 -143
rect 2323 -145 2325 -143
rect 40 -243 42 -241
rect 40 -250 42 -248
rect 80 -243 82 -241
rect 80 -250 82 -248
rect 90 -245 92 -243
rect 90 -252 92 -250
rect 168 -242 170 -240
rect 168 -249 170 -247
rect 180 -242 182 -240
rect 180 -249 182 -247
rect 258 -245 260 -243
rect 258 -252 260 -250
rect 299 -247 301 -245
rect 299 -254 301 -252
rect 347 -243 349 -241
rect 347 -250 349 -248
rect 357 -245 359 -243
rect 357 -252 359 -250
rect 435 -242 437 -240
rect 435 -249 437 -247
rect 447 -242 449 -240
rect 447 -249 449 -247
rect 525 -245 527 -243
rect 525 -252 527 -250
rect 566 -247 568 -245
rect 566 -254 568 -252
rect 614 -243 616 -241
rect 614 -250 616 -248
rect 624 -245 626 -243
rect 624 -252 626 -250
rect 702 -242 704 -240
rect 702 -249 704 -247
rect 714 -242 716 -240
rect 714 -249 716 -247
rect 792 -245 794 -243
rect 792 -252 794 -250
rect 833 -247 835 -245
rect 833 -254 835 -252
rect 881 -243 883 -241
rect 881 -250 883 -248
rect 891 -245 893 -243
rect 891 -252 893 -250
rect 969 -242 971 -240
rect 969 -249 971 -247
rect 981 -242 983 -240
rect 981 -249 983 -247
rect 1059 -245 1061 -243
rect 1059 -252 1061 -250
rect 1100 -247 1102 -245
rect 1100 -254 1102 -252
rect 1148 -243 1150 -241
rect 1148 -250 1150 -248
rect 1158 -245 1160 -243
rect 1158 -252 1160 -250
rect 1236 -242 1238 -240
rect 1236 -249 1238 -247
rect 1248 -242 1250 -240
rect 1248 -249 1250 -247
rect 1326 -245 1328 -243
rect 1326 -252 1328 -250
rect 1367 -247 1369 -245
rect 1367 -254 1369 -252
rect 1415 -243 1417 -241
rect 1415 -250 1417 -248
rect 1425 -245 1427 -243
rect 1425 -252 1427 -250
rect 1503 -242 1505 -240
rect 1503 -249 1505 -247
rect 1515 -242 1517 -240
rect 1515 -249 1517 -247
rect 1593 -245 1595 -243
rect 1593 -252 1595 -250
rect 1634 -247 1636 -245
rect 1634 -254 1636 -252
rect 1682 -243 1684 -241
rect 1682 -250 1684 -248
rect 1692 -245 1694 -243
rect 1692 -252 1694 -250
rect 1770 -242 1772 -240
rect 1770 -249 1772 -247
rect 1782 -242 1784 -240
rect 1782 -249 1784 -247
rect 1860 -245 1862 -243
rect 1860 -252 1862 -250
rect 1901 -247 1903 -245
rect 1901 -254 1903 -252
rect 1958 -250 1960 -248
rect 1978 -245 1980 -243
rect 1978 -252 1980 -250
rect 2056 -242 2058 -240
rect 2056 -249 2058 -247
rect 2068 -242 2070 -240
rect 2068 -249 2070 -247
rect 2146 -245 2148 -243
rect 2146 -252 2148 -250
rect 2187 -247 2189 -245
rect 2187 -254 2189 -252
rect 2255 -257 2257 -255
rect 2323 -257 2325 -255
<< alu0 >>
rect 8 289 14 296
rect 8 287 10 289
rect 12 287 14 289
rect 8 286 14 287
rect 19 289 23 291
rect 19 287 20 289
rect 22 287 23 289
rect 19 282 23 287
rect 28 287 34 296
rect 28 285 30 287
rect 32 285 34 287
rect 48 289 54 296
rect 48 287 50 289
rect 52 287 54 289
rect 48 286 54 287
rect 59 289 63 291
rect 59 287 60 289
rect 62 287 63 289
rect 28 284 34 285
rect 19 280 20 282
rect 22 281 23 282
rect 22 280 36 281
rect 19 277 36 280
rect 32 265 36 277
rect 32 263 33 265
rect 35 263 36 265
rect 32 258 36 263
rect 24 254 36 258
rect 59 282 63 287
rect 68 287 74 296
rect 99 294 101 296
rect 103 294 105 296
rect 99 293 105 294
rect 134 294 136 296
rect 138 294 140 296
rect 68 285 70 287
rect 72 285 74 287
rect 134 289 140 294
rect 156 294 158 296
rect 160 294 162 296
rect 134 287 136 289
rect 138 287 140 289
rect 134 286 140 287
rect 147 288 151 290
rect 147 286 148 288
rect 150 286 151 288
rect 156 289 162 294
rect 156 287 158 289
rect 160 287 162 289
rect 156 286 162 287
rect 188 294 190 296
rect 192 294 194 296
rect 188 289 194 294
rect 210 294 212 296
rect 214 294 216 296
rect 188 287 190 289
rect 192 287 194 289
rect 188 286 194 287
rect 199 288 203 290
rect 199 286 200 288
rect 202 286 203 288
rect 210 289 216 294
rect 245 294 247 296
rect 249 294 251 296
rect 245 293 251 294
rect 286 294 288 296
rect 290 294 292 296
rect 286 293 292 294
rect 210 287 212 289
rect 214 287 216 289
rect 210 286 216 287
rect 267 289 284 290
rect 267 287 269 289
rect 271 287 284 289
rect 267 286 284 287
rect 315 289 321 296
rect 315 287 317 289
rect 319 287 321 289
rect 315 286 321 287
rect 326 289 330 291
rect 326 287 327 289
rect 329 287 330 289
rect 68 284 74 285
rect 59 280 60 282
rect 62 281 63 282
rect 62 280 76 281
rect 59 277 76 280
rect 24 250 28 254
rect 39 251 40 253
rect 72 265 76 277
rect 72 263 73 265
rect 75 263 76 265
rect 72 258 76 263
rect 64 254 76 258
rect 8 249 28 250
rect 8 247 10 249
rect 12 247 28 249
rect 8 246 28 247
rect 64 250 68 254
rect 79 251 80 253
rect 48 249 68 250
rect 48 247 50 249
rect 52 247 68 249
rect 48 246 68 247
rect 104 282 128 286
rect 147 282 151 286
rect 102 278 108 282
rect 124 281 164 282
rect 124 279 148 281
rect 150 279 164 281
rect 102 268 106 278
rect 112 277 116 279
rect 124 278 164 279
rect 112 275 113 277
rect 115 275 116 277
rect 112 274 116 275
rect 102 266 103 268
rect 105 266 106 268
rect 102 264 106 266
rect 109 270 116 274
rect 109 259 113 270
rect 152 265 156 270
rect 152 263 153 265
rect 155 263 156 265
rect 95 258 113 259
rect 95 256 97 258
rect 99 257 113 258
rect 99 256 124 257
rect 95 255 120 256
rect 109 254 120 255
rect 122 254 124 256
rect 109 253 124 254
rect 129 256 133 258
rect 129 254 130 256
rect 132 254 133 256
rect 129 249 133 254
rect 152 261 156 263
rect 160 267 164 278
rect 160 265 166 267
rect 160 263 163 265
rect 165 263 166 265
rect 160 261 166 263
rect 160 258 164 261
rect 144 254 164 258
rect 144 250 148 254
rect 108 248 130 249
rect 99 245 103 247
rect 108 246 110 248
rect 112 247 130 248
rect 132 247 133 249
rect 112 246 133 247
rect 138 249 148 250
rect 138 247 140 249
rect 142 247 148 249
rect 138 246 148 247
rect 199 282 203 286
rect 222 282 246 286
rect 186 281 226 282
rect 186 279 200 281
rect 202 279 226 281
rect 186 278 226 279
rect 186 267 190 278
rect 234 277 238 279
rect 242 278 248 282
rect 234 275 235 277
rect 237 275 238 277
rect 234 274 238 275
rect 234 270 241 274
rect 184 265 190 267
rect 184 263 185 265
rect 187 263 190 265
rect 184 261 190 263
rect 194 265 198 270
rect 194 263 195 265
rect 197 263 198 265
rect 194 261 198 263
rect 186 258 190 261
rect 186 254 206 258
rect 202 250 206 254
rect 237 259 241 270
rect 244 268 248 278
rect 244 266 245 268
rect 247 266 248 268
rect 244 264 248 266
rect 237 258 255 259
rect 217 256 221 258
rect 237 257 251 258
rect 217 254 218 256
rect 220 254 221 256
rect 202 249 212 250
rect 202 247 208 249
rect 210 247 212 249
rect 202 246 212 247
rect 217 249 221 254
rect 226 256 251 257
rect 253 256 255 258
rect 226 254 228 256
rect 230 255 255 256
rect 230 254 241 255
rect 226 253 241 254
rect 280 282 284 286
rect 280 278 295 282
rect 270 269 276 270
rect 291 265 295 278
rect 298 275 299 286
rect 291 263 292 265
rect 294 263 295 265
rect 291 257 295 263
rect 326 282 330 287
rect 335 287 341 296
rect 366 294 368 296
rect 370 294 372 296
rect 366 293 372 294
rect 401 294 403 296
rect 405 294 407 296
rect 335 285 337 287
rect 339 285 341 287
rect 401 289 407 294
rect 423 294 425 296
rect 427 294 429 296
rect 401 287 403 289
rect 405 287 407 289
rect 401 286 407 287
rect 414 288 418 290
rect 414 286 415 288
rect 417 286 418 288
rect 423 289 429 294
rect 423 287 425 289
rect 427 287 429 289
rect 423 286 429 287
rect 455 294 457 296
rect 459 294 461 296
rect 455 289 461 294
rect 477 294 479 296
rect 481 294 483 296
rect 455 287 457 289
rect 459 287 461 289
rect 455 286 461 287
rect 466 288 470 290
rect 466 286 467 288
rect 469 286 470 288
rect 477 289 483 294
rect 512 294 514 296
rect 516 294 518 296
rect 512 293 518 294
rect 553 294 555 296
rect 557 294 559 296
rect 553 293 559 294
rect 477 287 479 289
rect 481 287 483 289
rect 477 286 483 287
rect 534 289 551 290
rect 534 287 536 289
rect 538 287 551 289
rect 534 286 551 287
rect 582 289 588 296
rect 582 287 584 289
rect 586 287 588 289
rect 582 286 588 287
rect 593 289 597 291
rect 593 287 594 289
rect 596 287 597 289
rect 335 284 341 285
rect 326 280 327 282
rect 329 281 330 282
rect 329 280 343 281
rect 326 277 343 280
rect 277 256 295 257
rect 277 254 279 256
rect 281 254 295 256
rect 277 253 295 254
rect 339 265 343 277
rect 339 263 340 265
rect 342 263 343 265
rect 339 258 343 263
rect 331 254 343 258
rect 331 250 335 254
rect 346 251 347 253
rect 217 247 218 249
rect 220 248 242 249
rect 220 247 238 248
rect 217 246 238 247
rect 240 246 242 248
rect 108 245 133 246
rect 217 245 242 246
rect 247 245 251 247
rect 315 249 335 250
rect 315 247 317 249
rect 319 247 335 249
rect 315 246 335 247
rect 371 282 395 286
rect 414 282 418 286
rect 369 278 375 282
rect 391 281 431 282
rect 391 279 415 281
rect 417 279 431 281
rect 369 268 373 278
rect 379 277 383 279
rect 391 278 431 279
rect 379 275 380 277
rect 382 275 383 277
rect 379 274 383 275
rect 369 266 370 268
rect 372 266 373 268
rect 369 264 373 266
rect 376 270 383 274
rect 376 259 380 270
rect 419 265 423 270
rect 419 263 420 265
rect 422 263 423 265
rect 362 258 380 259
rect 362 256 364 258
rect 366 257 380 258
rect 366 256 391 257
rect 362 255 387 256
rect 376 254 387 255
rect 389 254 391 256
rect 376 253 391 254
rect 396 256 400 258
rect 396 254 397 256
rect 399 254 400 256
rect 396 249 400 254
rect 419 261 423 263
rect 427 267 431 278
rect 427 265 433 267
rect 427 263 430 265
rect 432 263 433 265
rect 427 261 433 263
rect 427 258 431 261
rect 411 254 431 258
rect 411 250 415 254
rect 375 248 397 249
rect 366 245 370 247
rect 375 246 377 248
rect 379 247 397 248
rect 399 247 400 249
rect 379 246 400 247
rect 405 249 415 250
rect 405 247 407 249
rect 409 247 415 249
rect 405 246 415 247
rect 466 282 470 286
rect 489 282 513 286
rect 453 281 493 282
rect 453 279 467 281
rect 469 279 493 281
rect 453 278 493 279
rect 453 267 457 278
rect 501 277 505 279
rect 509 278 515 282
rect 501 275 502 277
rect 504 275 505 277
rect 501 274 505 275
rect 501 270 508 274
rect 451 265 457 267
rect 451 263 452 265
rect 454 263 457 265
rect 451 261 457 263
rect 461 265 465 270
rect 461 263 462 265
rect 464 263 465 265
rect 461 261 465 263
rect 453 258 457 261
rect 453 254 473 258
rect 469 250 473 254
rect 504 259 508 270
rect 511 268 515 278
rect 511 266 512 268
rect 514 266 515 268
rect 511 264 515 266
rect 504 258 522 259
rect 484 256 488 258
rect 504 257 518 258
rect 484 254 485 256
rect 487 254 488 256
rect 469 249 479 250
rect 469 247 475 249
rect 477 247 479 249
rect 469 246 479 247
rect 484 249 488 254
rect 493 256 518 257
rect 520 256 522 258
rect 493 254 495 256
rect 497 255 522 256
rect 497 254 508 255
rect 493 253 508 254
rect 547 282 551 286
rect 547 278 562 282
rect 537 269 543 270
rect 558 265 562 278
rect 565 275 566 286
rect 558 263 559 265
rect 561 263 562 265
rect 558 257 562 263
rect 593 282 597 287
rect 602 287 608 296
rect 633 294 635 296
rect 637 294 639 296
rect 633 293 639 294
rect 668 294 670 296
rect 672 294 674 296
rect 602 285 604 287
rect 606 285 608 287
rect 668 289 674 294
rect 690 294 692 296
rect 694 294 696 296
rect 668 287 670 289
rect 672 287 674 289
rect 668 286 674 287
rect 681 288 685 290
rect 681 286 682 288
rect 684 286 685 288
rect 690 289 696 294
rect 690 287 692 289
rect 694 287 696 289
rect 690 286 696 287
rect 722 294 724 296
rect 726 294 728 296
rect 722 289 728 294
rect 744 294 746 296
rect 748 294 750 296
rect 722 287 724 289
rect 726 287 728 289
rect 722 286 728 287
rect 733 288 737 290
rect 733 286 734 288
rect 736 286 737 288
rect 744 289 750 294
rect 779 294 781 296
rect 783 294 785 296
rect 779 293 785 294
rect 820 294 822 296
rect 824 294 826 296
rect 820 293 826 294
rect 744 287 746 289
rect 748 287 750 289
rect 744 286 750 287
rect 801 289 818 290
rect 801 287 803 289
rect 805 287 818 289
rect 801 286 818 287
rect 849 289 855 296
rect 849 287 851 289
rect 853 287 855 289
rect 849 286 855 287
rect 860 289 864 291
rect 860 287 861 289
rect 863 287 864 289
rect 602 284 608 285
rect 593 280 594 282
rect 596 281 597 282
rect 596 280 610 281
rect 593 277 610 280
rect 544 256 562 257
rect 544 254 546 256
rect 548 254 562 256
rect 544 253 562 254
rect 606 265 610 277
rect 606 263 607 265
rect 609 263 610 265
rect 606 258 610 263
rect 598 254 610 258
rect 598 250 602 254
rect 613 251 614 253
rect 484 247 485 249
rect 487 248 509 249
rect 487 247 505 248
rect 484 246 505 247
rect 507 246 509 248
rect 375 245 400 246
rect 484 245 509 246
rect 514 245 518 247
rect 582 249 602 250
rect 582 247 584 249
rect 586 247 602 249
rect 582 246 602 247
rect 638 282 662 286
rect 681 282 685 286
rect 636 278 642 282
rect 658 281 698 282
rect 658 279 682 281
rect 684 279 698 281
rect 636 268 640 278
rect 646 277 650 279
rect 658 278 698 279
rect 646 275 647 277
rect 649 275 650 277
rect 646 274 650 275
rect 636 266 637 268
rect 639 266 640 268
rect 636 264 640 266
rect 643 270 650 274
rect 643 259 647 270
rect 686 265 690 270
rect 686 263 687 265
rect 689 263 690 265
rect 629 258 647 259
rect 629 256 631 258
rect 633 257 647 258
rect 633 256 658 257
rect 629 255 654 256
rect 643 254 654 255
rect 656 254 658 256
rect 643 253 658 254
rect 663 256 667 258
rect 663 254 664 256
rect 666 254 667 256
rect 663 249 667 254
rect 686 261 690 263
rect 694 267 698 278
rect 694 265 700 267
rect 694 263 697 265
rect 699 263 700 265
rect 694 261 700 263
rect 694 258 698 261
rect 678 254 698 258
rect 678 250 682 254
rect 642 248 664 249
rect 633 245 637 247
rect 642 246 644 248
rect 646 247 664 248
rect 666 247 667 249
rect 646 246 667 247
rect 672 249 682 250
rect 672 247 674 249
rect 676 247 682 249
rect 672 246 682 247
rect 733 282 737 286
rect 756 282 780 286
rect 720 281 760 282
rect 720 279 734 281
rect 736 279 760 281
rect 720 278 760 279
rect 720 267 724 278
rect 768 277 772 279
rect 776 278 782 282
rect 768 275 769 277
rect 771 275 772 277
rect 768 274 772 275
rect 768 270 775 274
rect 718 265 724 267
rect 718 263 719 265
rect 721 263 724 265
rect 718 261 724 263
rect 728 265 732 270
rect 728 263 729 265
rect 731 263 732 265
rect 728 261 732 263
rect 720 258 724 261
rect 720 254 740 258
rect 736 250 740 254
rect 771 259 775 270
rect 778 268 782 278
rect 778 266 779 268
rect 781 266 782 268
rect 778 264 782 266
rect 771 258 789 259
rect 751 256 755 258
rect 771 257 785 258
rect 751 254 752 256
rect 754 254 755 256
rect 736 249 746 250
rect 736 247 742 249
rect 744 247 746 249
rect 736 246 746 247
rect 751 249 755 254
rect 760 256 785 257
rect 787 256 789 258
rect 760 254 762 256
rect 764 255 789 256
rect 814 282 818 286
rect 814 278 829 282
rect 804 269 810 270
rect 764 254 775 255
rect 760 253 775 254
rect 825 265 829 278
rect 832 275 833 286
rect 825 263 826 265
rect 828 263 829 265
rect 825 257 829 263
rect 860 282 864 287
rect 869 287 875 296
rect 900 294 902 296
rect 904 294 906 296
rect 900 293 906 294
rect 935 294 937 296
rect 939 294 941 296
rect 869 285 871 287
rect 873 285 875 287
rect 935 289 941 294
rect 957 294 959 296
rect 961 294 963 296
rect 935 287 937 289
rect 939 287 941 289
rect 935 286 941 287
rect 948 288 952 290
rect 948 286 949 288
rect 951 286 952 288
rect 957 289 963 294
rect 957 287 959 289
rect 961 287 963 289
rect 957 286 963 287
rect 989 294 991 296
rect 993 294 995 296
rect 989 289 995 294
rect 1011 294 1013 296
rect 1015 294 1017 296
rect 989 287 991 289
rect 993 287 995 289
rect 989 286 995 287
rect 1000 288 1004 290
rect 1000 286 1001 288
rect 1003 286 1004 288
rect 1011 289 1017 294
rect 1046 294 1048 296
rect 1050 294 1052 296
rect 1046 293 1052 294
rect 1087 294 1089 296
rect 1091 294 1093 296
rect 1087 293 1093 294
rect 1011 287 1013 289
rect 1015 287 1017 289
rect 1011 286 1017 287
rect 1068 289 1085 290
rect 1068 287 1070 289
rect 1072 287 1085 289
rect 1068 286 1085 287
rect 1116 289 1122 296
rect 1116 287 1118 289
rect 1120 287 1122 289
rect 1116 286 1122 287
rect 1127 289 1131 291
rect 1127 287 1128 289
rect 1130 287 1131 289
rect 869 284 875 285
rect 860 280 861 282
rect 863 281 864 282
rect 863 280 877 281
rect 860 277 877 280
rect 811 256 829 257
rect 811 254 813 256
rect 815 254 829 256
rect 811 253 829 254
rect 873 265 877 277
rect 873 263 874 265
rect 876 263 877 265
rect 873 258 877 263
rect 865 254 877 258
rect 865 250 869 254
rect 880 251 881 253
rect 751 247 752 249
rect 754 248 776 249
rect 754 247 772 248
rect 751 246 772 247
rect 774 246 776 248
rect 642 245 667 246
rect 751 245 776 246
rect 781 245 785 247
rect 849 249 869 250
rect 849 247 851 249
rect 853 247 869 249
rect 849 246 869 247
rect 905 282 929 286
rect 948 282 952 286
rect 903 278 909 282
rect 925 281 965 282
rect 925 279 949 281
rect 951 279 965 281
rect 903 268 907 278
rect 913 277 917 279
rect 925 278 965 279
rect 913 275 914 277
rect 916 275 917 277
rect 913 274 917 275
rect 903 266 904 268
rect 906 266 907 268
rect 903 264 907 266
rect 910 270 917 274
rect 910 259 914 270
rect 953 265 957 270
rect 953 263 954 265
rect 956 263 957 265
rect 896 258 914 259
rect 896 256 898 258
rect 900 257 914 258
rect 900 256 925 257
rect 896 255 921 256
rect 910 254 921 255
rect 923 254 925 256
rect 910 253 925 254
rect 930 256 934 258
rect 930 254 931 256
rect 933 254 934 256
rect 930 249 934 254
rect 953 261 957 263
rect 961 267 965 278
rect 961 265 967 267
rect 961 263 964 265
rect 966 263 967 265
rect 961 261 967 263
rect 961 258 965 261
rect 945 254 965 258
rect 945 250 949 254
rect 909 248 931 249
rect 900 245 904 247
rect 909 246 911 248
rect 913 247 931 248
rect 933 247 934 249
rect 913 246 934 247
rect 939 249 949 250
rect 939 247 941 249
rect 943 247 949 249
rect 939 246 949 247
rect 1000 282 1004 286
rect 1023 282 1047 286
rect 987 281 1027 282
rect 987 279 1001 281
rect 1003 279 1027 281
rect 987 278 1027 279
rect 987 267 991 278
rect 1035 277 1039 279
rect 1043 278 1049 282
rect 1035 275 1036 277
rect 1038 275 1039 277
rect 1035 274 1039 275
rect 1035 270 1042 274
rect 985 265 991 267
rect 985 263 986 265
rect 988 263 991 265
rect 985 261 991 263
rect 995 265 999 270
rect 995 263 996 265
rect 998 263 999 265
rect 995 261 999 263
rect 987 258 991 261
rect 987 254 1007 258
rect 1003 250 1007 254
rect 1038 259 1042 270
rect 1045 268 1049 278
rect 1045 266 1046 268
rect 1048 266 1049 268
rect 1045 264 1049 266
rect 1038 258 1056 259
rect 1018 256 1022 258
rect 1038 257 1052 258
rect 1018 254 1019 256
rect 1021 254 1022 256
rect 1003 249 1013 250
rect 1003 247 1009 249
rect 1011 247 1013 249
rect 1003 246 1013 247
rect 1018 249 1022 254
rect 1027 256 1052 257
rect 1054 256 1056 258
rect 1027 254 1029 256
rect 1031 255 1056 256
rect 1081 282 1085 286
rect 1081 278 1096 282
rect 1071 269 1077 270
rect 1031 254 1042 255
rect 1027 253 1042 254
rect 1092 265 1096 278
rect 1099 275 1100 286
rect 1092 263 1093 265
rect 1095 263 1096 265
rect 1092 257 1096 263
rect 1127 282 1131 287
rect 1136 287 1142 296
rect 1167 294 1169 296
rect 1171 294 1173 296
rect 1167 293 1173 294
rect 1202 294 1204 296
rect 1206 294 1208 296
rect 1136 285 1138 287
rect 1140 285 1142 287
rect 1202 289 1208 294
rect 1224 294 1226 296
rect 1228 294 1230 296
rect 1202 287 1204 289
rect 1206 287 1208 289
rect 1202 286 1208 287
rect 1215 288 1219 290
rect 1215 286 1216 288
rect 1218 286 1219 288
rect 1224 289 1230 294
rect 1224 287 1226 289
rect 1228 287 1230 289
rect 1224 286 1230 287
rect 1256 294 1258 296
rect 1260 294 1262 296
rect 1256 289 1262 294
rect 1278 294 1280 296
rect 1282 294 1284 296
rect 1256 287 1258 289
rect 1260 287 1262 289
rect 1256 286 1262 287
rect 1267 288 1271 290
rect 1267 286 1268 288
rect 1270 286 1271 288
rect 1278 289 1284 294
rect 1313 294 1315 296
rect 1317 294 1319 296
rect 1313 293 1319 294
rect 1354 294 1356 296
rect 1358 294 1360 296
rect 1354 293 1360 294
rect 1278 287 1280 289
rect 1282 287 1284 289
rect 1278 286 1284 287
rect 1335 289 1352 290
rect 1335 287 1337 289
rect 1339 287 1352 289
rect 1335 286 1352 287
rect 1383 289 1389 296
rect 1383 287 1385 289
rect 1387 287 1389 289
rect 1383 286 1389 287
rect 1394 289 1398 291
rect 1394 287 1395 289
rect 1397 287 1398 289
rect 1136 284 1142 285
rect 1127 280 1128 282
rect 1130 281 1131 282
rect 1130 280 1144 281
rect 1127 277 1144 280
rect 1078 256 1096 257
rect 1078 254 1080 256
rect 1082 254 1096 256
rect 1078 253 1096 254
rect 1140 265 1144 277
rect 1140 263 1141 265
rect 1143 263 1144 265
rect 1140 258 1144 263
rect 1132 254 1144 258
rect 1132 250 1136 254
rect 1147 251 1148 253
rect 1018 247 1019 249
rect 1021 248 1043 249
rect 1021 247 1039 248
rect 1018 246 1039 247
rect 1041 246 1043 248
rect 909 245 934 246
rect 1018 245 1043 246
rect 1048 245 1052 247
rect 1116 249 1136 250
rect 1116 247 1118 249
rect 1120 247 1136 249
rect 1116 246 1136 247
rect 1172 282 1196 286
rect 1215 282 1219 286
rect 1170 278 1176 282
rect 1192 281 1232 282
rect 1192 279 1216 281
rect 1218 279 1232 281
rect 1170 268 1174 278
rect 1180 277 1184 279
rect 1192 278 1232 279
rect 1180 275 1181 277
rect 1183 275 1184 277
rect 1180 274 1184 275
rect 1170 266 1171 268
rect 1173 266 1174 268
rect 1170 264 1174 266
rect 1177 270 1184 274
rect 1177 259 1181 270
rect 1220 265 1224 270
rect 1220 263 1221 265
rect 1223 263 1224 265
rect 1163 258 1181 259
rect 1163 256 1165 258
rect 1167 257 1181 258
rect 1167 256 1192 257
rect 1163 255 1188 256
rect 1177 254 1188 255
rect 1190 254 1192 256
rect 1177 253 1192 254
rect 1197 256 1201 258
rect 1197 254 1198 256
rect 1200 254 1201 256
rect 1197 249 1201 254
rect 1220 261 1224 263
rect 1228 267 1232 278
rect 1228 265 1234 267
rect 1228 263 1231 265
rect 1233 263 1234 265
rect 1228 261 1234 263
rect 1228 258 1232 261
rect 1212 254 1232 258
rect 1212 250 1216 254
rect 1176 248 1198 249
rect 1167 245 1171 247
rect 1176 246 1178 248
rect 1180 247 1198 248
rect 1200 247 1201 249
rect 1180 246 1201 247
rect 1206 249 1216 250
rect 1206 247 1208 249
rect 1210 247 1216 249
rect 1206 246 1216 247
rect 1267 282 1271 286
rect 1290 282 1314 286
rect 1254 281 1294 282
rect 1254 279 1268 281
rect 1270 279 1294 281
rect 1254 278 1294 279
rect 1254 267 1258 278
rect 1302 277 1306 279
rect 1310 278 1316 282
rect 1302 275 1303 277
rect 1305 275 1306 277
rect 1302 274 1306 275
rect 1302 270 1309 274
rect 1252 265 1258 267
rect 1252 263 1253 265
rect 1255 263 1258 265
rect 1252 261 1258 263
rect 1262 265 1266 270
rect 1262 263 1263 265
rect 1265 263 1266 265
rect 1262 261 1266 263
rect 1254 258 1258 261
rect 1254 254 1274 258
rect 1270 250 1274 254
rect 1305 259 1309 270
rect 1312 268 1316 278
rect 1312 266 1313 268
rect 1315 266 1316 268
rect 1312 264 1316 266
rect 1305 258 1323 259
rect 1285 256 1289 258
rect 1305 257 1319 258
rect 1285 254 1286 256
rect 1288 254 1289 256
rect 1270 249 1280 250
rect 1270 247 1276 249
rect 1278 247 1280 249
rect 1270 246 1280 247
rect 1285 249 1289 254
rect 1294 256 1319 257
rect 1321 256 1323 258
rect 1294 254 1296 256
rect 1298 255 1323 256
rect 1298 254 1309 255
rect 1294 253 1309 254
rect 1348 282 1352 286
rect 1348 278 1363 282
rect 1338 269 1344 270
rect 1359 265 1363 278
rect 1366 275 1367 286
rect 1359 263 1360 265
rect 1362 263 1363 265
rect 1359 257 1363 263
rect 1394 282 1398 287
rect 1403 287 1409 296
rect 1434 294 1436 296
rect 1438 294 1440 296
rect 1434 293 1440 294
rect 1469 294 1471 296
rect 1473 294 1475 296
rect 1403 285 1405 287
rect 1407 285 1409 287
rect 1469 289 1475 294
rect 1491 294 1493 296
rect 1495 294 1497 296
rect 1469 287 1471 289
rect 1473 287 1475 289
rect 1469 286 1475 287
rect 1482 288 1486 290
rect 1482 286 1483 288
rect 1485 286 1486 288
rect 1491 289 1497 294
rect 1491 287 1493 289
rect 1495 287 1497 289
rect 1491 286 1497 287
rect 1523 294 1525 296
rect 1527 294 1529 296
rect 1523 289 1529 294
rect 1545 294 1547 296
rect 1549 294 1551 296
rect 1523 287 1525 289
rect 1527 287 1529 289
rect 1523 286 1529 287
rect 1534 288 1538 290
rect 1534 286 1535 288
rect 1537 286 1538 288
rect 1545 289 1551 294
rect 1580 294 1582 296
rect 1584 294 1586 296
rect 1580 293 1586 294
rect 1621 294 1623 296
rect 1625 294 1627 296
rect 1621 293 1627 294
rect 1545 287 1547 289
rect 1549 287 1551 289
rect 1545 286 1551 287
rect 1602 289 1619 290
rect 1602 287 1604 289
rect 1606 287 1619 289
rect 1602 286 1619 287
rect 1650 289 1656 296
rect 1650 287 1652 289
rect 1654 287 1656 289
rect 1650 286 1656 287
rect 1661 289 1665 291
rect 1661 287 1662 289
rect 1664 287 1665 289
rect 1403 284 1409 285
rect 1394 280 1395 282
rect 1397 281 1398 282
rect 1397 280 1411 281
rect 1394 277 1411 280
rect 1345 256 1363 257
rect 1345 254 1347 256
rect 1349 254 1363 256
rect 1345 253 1363 254
rect 1407 265 1411 277
rect 1407 263 1408 265
rect 1410 263 1411 265
rect 1407 258 1411 263
rect 1399 254 1411 258
rect 1399 250 1403 254
rect 1414 251 1415 253
rect 1285 247 1286 249
rect 1288 248 1310 249
rect 1288 247 1306 248
rect 1285 246 1306 247
rect 1308 246 1310 248
rect 1176 245 1201 246
rect 1285 245 1310 246
rect 1315 245 1319 247
rect 1383 249 1403 250
rect 1383 247 1385 249
rect 1387 247 1403 249
rect 1383 246 1403 247
rect 1439 282 1463 286
rect 1482 282 1486 286
rect 1437 278 1443 282
rect 1459 281 1499 282
rect 1459 279 1483 281
rect 1485 279 1499 281
rect 1437 268 1441 278
rect 1447 277 1451 279
rect 1459 278 1499 279
rect 1447 275 1448 277
rect 1450 275 1451 277
rect 1447 274 1451 275
rect 1437 266 1438 268
rect 1440 266 1441 268
rect 1437 264 1441 266
rect 1444 270 1451 274
rect 1444 259 1448 270
rect 1487 265 1491 270
rect 1487 263 1488 265
rect 1490 263 1491 265
rect 1430 258 1448 259
rect 1430 256 1432 258
rect 1434 257 1448 258
rect 1434 256 1459 257
rect 1430 255 1455 256
rect 1444 254 1455 255
rect 1457 254 1459 256
rect 1444 253 1459 254
rect 1464 256 1468 258
rect 1464 254 1465 256
rect 1467 254 1468 256
rect 1464 249 1468 254
rect 1487 261 1491 263
rect 1495 267 1499 278
rect 1495 265 1501 267
rect 1495 263 1498 265
rect 1500 263 1501 265
rect 1495 261 1501 263
rect 1495 258 1499 261
rect 1479 254 1499 258
rect 1479 250 1483 254
rect 1443 248 1465 249
rect 1434 245 1438 247
rect 1443 246 1445 248
rect 1447 247 1465 248
rect 1467 247 1468 249
rect 1447 246 1468 247
rect 1473 249 1483 250
rect 1473 247 1475 249
rect 1477 247 1483 249
rect 1473 246 1483 247
rect 1534 282 1538 286
rect 1557 282 1581 286
rect 1521 281 1561 282
rect 1521 279 1535 281
rect 1537 279 1561 281
rect 1521 278 1561 279
rect 1521 267 1525 278
rect 1569 277 1573 279
rect 1577 278 1583 282
rect 1569 275 1570 277
rect 1572 275 1573 277
rect 1569 274 1573 275
rect 1569 270 1576 274
rect 1519 265 1525 267
rect 1519 263 1520 265
rect 1522 263 1525 265
rect 1519 261 1525 263
rect 1529 265 1533 270
rect 1529 263 1530 265
rect 1532 263 1533 265
rect 1529 261 1533 263
rect 1521 258 1525 261
rect 1521 254 1541 258
rect 1537 250 1541 254
rect 1572 259 1576 270
rect 1579 268 1583 278
rect 1579 266 1580 268
rect 1582 266 1583 268
rect 1579 264 1583 266
rect 1572 258 1590 259
rect 1552 256 1556 258
rect 1572 257 1586 258
rect 1552 254 1553 256
rect 1555 254 1556 256
rect 1537 249 1547 250
rect 1537 247 1543 249
rect 1545 247 1547 249
rect 1537 246 1547 247
rect 1552 249 1556 254
rect 1561 256 1586 257
rect 1588 256 1590 258
rect 1561 254 1563 256
rect 1565 255 1590 256
rect 1565 254 1576 255
rect 1561 253 1576 254
rect 1615 282 1619 286
rect 1615 278 1630 282
rect 1605 269 1611 270
rect 1626 265 1630 278
rect 1633 275 1634 286
rect 1626 263 1627 265
rect 1629 263 1630 265
rect 1626 257 1630 263
rect 1661 282 1665 287
rect 1670 287 1676 296
rect 1701 294 1703 296
rect 1705 294 1707 296
rect 1701 293 1707 294
rect 1736 294 1738 296
rect 1740 294 1742 296
rect 1670 285 1672 287
rect 1674 285 1676 287
rect 1736 289 1742 294
rect 1758 294 1760 296
rect 1762 294 1764 296
rect 1736 287 1738 289
rect 1740 287 1742 289
rect 1736 286 1742 287
rect 1749 288 1753 290
rect 1749 286 1750 288
rect 1752 286 1753 288
rect 1758 289 1764 294
rect 1758 287 1760 289
rect 1762 287 1764 289
rect 1758 286 1764 287
rect 1790 294 1792 296
rect 1794 294 1796 296
rect 1790 289 1796 294
rect 1812 294 1814 296
rect 1816 294 1818 296
rect 1790 287 1792 289
rect 1794 287 1796 289
rect 1790 286 1796 287
rect 1801 288 1805 290
rect 1801 286 1802 288
rect 1804 286 1805 288
rect 1812 289 1818 294
rect 1847 294 1849 296
rect 1851 294 1853 296
rect 1847 293 1853 294
rect 1888 294 1890 296
rect 1892 294 1894 296
rect 1888 293 1894 294
rect 1931 294 1932 296
rect 1934 294 1935 296
rect 1812 287 1814 289
rect 1816 287 1818 289
rect 1812 286 1818 287
rect 1869 289 1886 290
rect 1869 287 1871 289
rect 1873 287 1886 289
rect 1869 286 1886 287
rect 1670 284 1676 285
rect 1661 280 1662 282
rect 1664 281 1665 282
rect 1664 280 1678 281
rect 1661 277 1678 280
rect 1612 256 1630 257
rect 1612 254 1614 256
rect 1616 254 1630 256
rect 1612 253 1630 254
rect 1674 265 1678 277
rect 1674 263 1675 265
rect 1677 263 1678 265
rect 1674 258 1678 263
rect 1666 254 1678 258
rect 1666 250 1670 254
rect 1681 251 1682 253
rect 1552 247 1553 249
rect 1555 248 1577 249
rect 1555 247 1573 248
rect 1552 246 1573 247
rect 1575 246 1577 248
rect 1443 245 1468 246
rect 1552 245 1577 246
rect 1582 245 1586 247
rect 1650 249 1670 250
rect 1650 247 1652 249
rect 1654 247 1670 249
rect 1650 246 1670 247
rect 1706 282 1730 286
rect 1749 282 1753 286
rect 1704 278 1710 282
rect 1726 281 1766 282
rect 1726 279 1750 281
rect 1752 279 1766 281
rect 1704 268 1708 278
rect 1714 277 1718 279
rect 1726 278 1766 279
rect 1714 275 1715 277
rect 1717 275 1718 277
rect 1714 274 1718 275
rect 1704 266 1705 268
rect 1707 266 1708 268
rect 1704 264 1708 266
rect 1711 270 1718 274
rect 1711 259 1715 270
rect 1754 265 1758 270
rect 1754 263 1755 265
rect 1757 263 1758 265
rect 1697 258 1715 259
rect 1697 256 1699 258
rect 1701 257 1715 258
rect 1701 256 1726 257
rect 1697 255 1722 256
rect 1711 254 1722 255
rect 1724 254 1726 256
rect 1711 253 1726 254
rect 1731 256 1735 258
rect 1731 254 1732 256
rect 1734 254 1735 256
rect 1731 249 1735 254
rect 1754 261 1758 263
rect 1762 267 1766 278
rect 1762 265 1768 267
rect 1762 263 1765 265
rect 1767 263 1768 265
rect 1762 261 1768 263
rect 1762 258 1766 261
rect 1746 254 1766 258
rect 1746 250 1750 254
rect 1710 248 1732 249
rect 1701 245 1705 247
rect 1710 246 1712 248
rect 1714 247 1732 248
rect 1734 247 1735 249
rect 1714 246 1735 247
rect 1740 249 1750 250
rect 1740 247 1742 249
rect 1744 247 1750 249
rect 1740 246 1750 247
rect 1801 282 1805 286
rect 1824 282 1848 286
rect 1788 281 1828 282
rect 1788 279 1802 281
rect 1804 279 1828 281
rect 1788 278 1828 279
rect 1788 267 1792 278
rect 1836 277 1840 279
rect 1844 278 1850 282
rect 1836 275 1837 277
rect 1839 275 1840 277
rect 1836 274 1840 275
rect 1836 270 1843 274
rect 1786 265 1792 267
rect 1786 263 1787 265
rect 1789 263 1792 265
rect 1786 261 1792 263
rect 1796 265 1800 270
rect 1796 263 1797 265
rect 1799 263 1800 265
rect 1796 261 1800 263
rect 1788 258 1792 261
rect 1788 254 1808 258
rect 1804 250 1808 254
rect 1839 259 1843 270
rect 1846 268 1850 278
rect 1846 266 1847 268
rect 1849 266 1850 268
rect 1846 264 1850 266
rect 1839 258 1857 259
rect 1819 256 1823 258
rect 1839 257 1853 258
rect 1819 254 1820 256
rect 1822 254 1823 256
rect 1804 249 1814 250
rect 1804 247 1810 249
rect 1812 247 1814 249
rect 1804 246 1814 247
rect 1819 249 1823 254
rect 1828 256 1853 257
rect 1855 256 1857 258
rect 1828 254 1830 256
rect 1832 255 1857 256
rect 1832 254 1843 255
rect 1828 253 1843 254
rect 1882 282 1886 286
rect 1882 278 1897 282
rect 1872 269 1878 270
rect 1893 265 1897 278
rect 1900 275 1901 286
rect 1893 263 1894 265
rect 1896 263 1897 265
rect 1893 257 1897 263
rect 1931 289 1935 294
rect 1987 294 1989 296
rect 1991 294 1993 296
rect 1987 293 1993 294
rect 2022 294 2024 296
rect 2026 294 2028 296
rect 1931 287 1932 289
rect 1934 287 1935 289
rect 1931 285 1935 287
rect 1939 290 1972 291
rect 1939 288 1968 290
rect 1970 288 1972 290
rect 1939 287 1972 288
rect 2022 289 2028 294
rect 2044 294 2046 296
rect 2048 294 2050 296
rect 2022 287 2024 289
rect 2026 287 2028 289
rect 1939 276 1943 287
rect 2022 286 2028 287
rect 2035 288 2039 290
rect 2035 286 2036 288
rect 2038 286 2039 288
rect 2044 289 2050 294
rect 2044 287 2046 289
rect 2048 287 2050 289
rect 2044 286 2050 287
rect 2076 294 2078 296
rect 2080 294 2082 296
rect 2076 289 2082 294
rect 2098 294 2100 296
rect 2102 294 2104 296
rect 2076 287 2078 289
rect 2080 287 2082 289
rect 2076 286 2082 287
rect 2087 288 2091 290
rect 2087 286 2088 288
rect 2090 286 2091 288
rect 2098 289 2104 294
rect 2133 294 2135 296
rect 2137 294 2139 296
rect 2133 293 2139 294
rect 2174 294 2176 296
rect 2178 294 2180 296
rect 2174 293 2180 294
rect 2210 294 2211 296
rect 2213 294 2214 296
rect 2210 292 2214 294
rect 2243 294 2245 296
rect 2247 294 2249 296
rect 2243 293 2249 294
rect 2278 294 2279 296
rect 2281 294 2282 296
rect 2278 292 2282 294
rect 2311 294 2313 296
rect 2315 294 2317 296
rect 2311 293 2317 294
rect 2098 287 2100 289
rect 2102 287 2104 289
rect 2098 286 2104 287
rect 2155 289 2172 290
rect 2155 287 2157 289
rect 2159 287 2172 289
rect 2155 286 2172 287
rect 1920 275 1943 276
rect 1920 273 1922 275
rect 1924 273 1943 275
rect 1920 272 1943 273
rect 1920 266 1924 272
rect 1879 256 1897 257
rect 1879 254 1881 256
rect 1883 254 1897 256
rect 1879 253 1897 254
rect 1913 262 1924 266
rect 1913 256 1917 262
rect 1939 266 1943 272
rect 1947 282 1951 284
rect 1947 280 1948 282
rect 1950 280 1951 282
rect 1947 275 1951 280
rect 1947 273 1948 275
rect 1950 274 1951 275
rect 1950 273 1963 274
rect 1947 270 1963 273
rect 1959 268 1963 270
rect 1959 266 1964 268
rect 1939 265 1955 266
rect 1939 263 1951 265
rect 1953 263 1955 265
rect 1939 262 1955 263
rect 1959 264 1961 266
rect 1963 264 1964 266
rect 1959 262 1964 264
rect 1913 254 1914 256
rect 1916 254 1917 256
rect 1913 252 1917 254
rect 1959 258 1963 262
rect 1939 254 1963 258
rect 1939 251 1943 254
rect 1939 249 1940 251
rect 1942 249 1943 251
rect 1819 247 1820 249
rect 1822 248 1844 249
rect 1822 247 1840 248
rect 1819 246 1840 247
rect 1842 246 1844 248
rect 1710 245 1735 246
rect 1819 245 1844 246
rect 1849 245 1853 247
rect 1926 248 1932 249
rect 1926 246 1928 248
rect 1930 246 1932 248
rect 1939 247 1943 249
rect 1992 282 2016 286
rect 2035 282 2039 286
rect 1990 278 1996 282
rect 2012 281 2052 282
rect 2012 279 2036 281
rect 2038 279 2052 281
rect 1990 268 1994 278
rect 2000 277 2004 279
rect 2012 278 2052 279
rect 2000 275 2001 277
rect 2003 275 2004 277
rect 2000 274 2004 275
rect 1990 266 1991 268
rect 1993 266 1994 268
rect 1990 264 1994 266
rect 1997 270 2004 274
rect 1997 259 2001 270
rect 2040 265 2044 270
rect 2040 263 2041 265
rect 2043 263 2044 265
rect 1983 258 2001 259
rect 1983 256 1985 258
rect 1987 257 2001 258
rect 1987 256 2012 257
rect 1983 255 2008 256
rect 1997 254 2008 255
rect 2010 254 2012 256
rect 1997 253 2012 254
rect 2017 256 2021 258
rect 2017 254 2018 256
rect 2020 254 2021 256
rect 2017 249 2021 254
rect 2040 261 2044 263
rect 2048 267 2052 278
rect 2048 265 2054 267
rect 2048 263 2051 265
rect 2053 263 2054 265
rect 2048 261 2054 263
rect 2048 258 2052 261
rect 2032 254 2052 258
rect 2032 250 2036 254
rect 1996 248 2018 249
rect 99 243 100 245
rect 102 243 103 245
rect 247 243 248 245
rect 250 243 251 245
rect 99 240 103 243
rect 155 242 161 243
rect 155 240 157 242
rect 159 240 161 242
rect 189 242 195 243
rect 189 240 191 242
rect 193 240 195 242
rect 247 240 251 243
rect 267 243 273 244
rect 267 241 269 243
rect 271 241 273 243
rect 267 240 273 241
rect 286 243 292 244
rect 286 241 288 243
rect 290 241 292 243
rect 286 240 292 241
rect 366 243 367 245
rect 369 243 370 245
rect 514 243 515 245
rect 517 243 518 245
rect 366 240 370 243
rect 422 242 428 243
rect 422 240 424 242
rect 426 240 428 242
rect 456 242 462 243
rect 456 240 458 242
rect 460 240 462 242
rect 514 240 518 243
rect 534 243 540 244
rect 534 241 536 243
rect 538 241 540 243
rect 534 240 540 241
rect 553 243 559 244
rect 553 241 555 243
rect 557 241 559 243
rect 553 240 559 241
rect 633 243 634 245
rect 636 243 637 245
rect 781 243 782 245
rect 784 243 785 245
rect 633 240 637 243
rect 689 242 695 243
rect 689 240 691 242
rect 693 240 695 242
rect 723 242 729 243
rect 723 240 725 242
rect 727 240 729 242
rect 781 240 785 243
rect 801 243 807 244
rect 801 241 803 243
rect 805 241 807 243
rect 801 240 807 241
rect 820 243 826 244
rect 820 241 822 243
rect 824 241 826 243
rect 820 240 826 241
rect 900 243 901 245
rect 903 243 904 245
rect 1048 243 1049 245
rect 1051 243 1052 245
rect 900 240 904 243
rect 956 242 962 243
rect 956 240 958 242
rect 960 240 962 242
rect 990 242 996 243
rect 990 240 992 242
rect 994 240 996 242
rect 1048 240 1052 243
rect 1068 243 1074 244
rect 1068 241 1070 243
rect 1072 241 1074 243
rect 1068 240 1074 241
rect 1087 243 1093 244
rect 1087 241 1089 243
rect 1091 241 1093 243
rect 1087 240 1093 241
rect 1167 243 1168 245
rect 1170 243 1171 245
rect 1315 243 1316 245
rect 1318 243 1319 245
rect 1167 240 1171 243
rect 1223 242 1229 243
rect 1223 240 1225 242
rect 1227 240 1229 242
rect 1257 242 1263 243
rect 1257 240 1259 242
rect 1261 240 1263 242
rect 1315 240 1319 243
rect 1335 243 1341 244
rect 1335 241 1337 243
rect 1339 241 1341 243
rect 1335 240 1341 241
rect 1354 243 1360 244
rect 1354 241 1356 243
rect 1358 241 1360 243
rect 1354 240 1360 241
rect 1434 243 1435 245
rect 1437 243 1438 245
rect 1582 243 1583 245
rect 1585 243 1586 245
rect 1434 240 1438 243
rect 1490 242 1496 243
rect 1490 240 1492 242
rect 1494 240 1496 242
rect 1524 242 1530 243
rect 1524 240 1526 242
rect 1528 240 1530 242
rect 1582 240 1586 243
rect 1602 243 1608 244
rect 1602 241 1604 243
rect 1606 241 1608 243
rect 1602 240 1608 241
rect 1621 243 1627 244
rect 1621 241 1623 243
rect 1625 241 1627 243
rect 1621 240 1627 241
rect 1701 243 1702 245
rect 1704 243 1705 245
rect 1849 243 1850 245
rect 1852 243 1853 245
rect 1701 240 1705 243
rect 1757 242 1763 243
rect 1757 240 1759 242
rect 1761 240 1763 242
rect 1791 242 1797 243
rect 1791 240 1793 242
rect 1795 240 1797 242
rect 1849 240 1853 243
rect 1869 243 1875 244
rect 1869 241 1871 243
rect 1873 241 1875 243
rect 1869 240 1875 241
rect 1888 243 1894 244
rect 1888 241 1890 243
rect 1892 241 1894 243
rect 1888 240 1894 241
rect 1926 240 1932 246
rect 1987 245 1991 247
rect 1996 246 1998 248
rect 2000 247 2018 248
rect 2020 247 2021 249
rect 2000 246 2021 247
rect 2026 249 2036 250
rect 2026 247 2028 249
rect 2030 247 2036 249
rect 2026 246 2036 247
rect 2087 282 2091 286
rect 2110 282 2134 286
rect 2074 281 2114 282
rect 2074 279 2088 281
rect 2090 279 2114 281
rect 2074 278 2114 279
rect 2074 267 2078 278
rect 2122 277 2126 279
rect 2130 278 2136 282
rect 2122 275 2123 277
rect 2125 275 2126 277
rect 2122 274 2126 275
rect 2122 270 2129 274
rect 2072 265 2078 267
rect 2072 263 2073 265
rect 2075 263 2078 265
rect 2072 261 2078 263
rect 2082 265 2086 270
rect 2082 263 2083 265
rect 2085 263 2086 265
rect 2082 261 2086 263
rect 2074 258 2078 261
rect 2074 254 2094 258
rect 2090 250 2094 254
rect 2125 259 2129 270
rect 2132 268 2136 278
rect 2132 266 2133 268
rect 2135 266 2136 268
rect 2132 264 2136 266
rect 2125 258 2143 259
rect 2105 256 2109 258
rect 2125 257 2139 258
rect 2105 254 2106 256
rect 2108 254 2109 256
rect 2090 249 2100 250
rect 2090 247 2096 249
rect 2098 247 2100 249
rect 2090 246 2100 247
rect 2105 249 2109 254
rect 2114 256 2139 257
rect 2141 256 2143 258
rect 2114 254 2116 256
rect 2118 255 2143 256
rect 2168 282 2172 286
rect 2168 278 2183 282
rect 2158 269 2164 270
rect 2118 254 2129 255
rect 2114 253 2129 254
rect 2179 265 2183 278
rect 2186 275 2187 286
rect 2226 286 2239 287
rect 2226 284 2228 286
rect 2230 284 2239 286
rect 2226 283 2239 284
rect 2235 279 2251 283
rect 2179 263 2180 265
rect 2182 263 2183 265
rect 2179 257 2183 263
rect 2223 275 2227 277
rect 2165 256 2183 257
rect 2165 254 2167 256
rect 2169 254 2183 256
rect 2165 253 2183 254
rect 2199 274 2224 275
rect 2199 272 2201 274
rect 2203 273 2224 274
rect 2226 273 2227 275
rect 2203 272 2227 273
rect 2199 271 2227 272
rect 2105 247 2106 249
rect 2108 248 2130 249
rect 2108 247 2126 248
rect 2105 246 2126 247
rect 2128 246 2130 248
rect 2199 251 2203 271
rect 2223 261 2227 271
rect 2243 266 2244 272
rect 2247 262 2251 279
rect 2223 259 2234 261
rect 2223 257 2231 259
rect 2233 257 2234 259
rect 2247 260 2252 262
rect 2247 258 2249 260
rect 2251 258 2252 260
rect 2223 255 2234 257
rect 2237 256 2252 258
rect 2237 254 2251 256
rect 2199 250 2205 251
rect 2199 248 2201 250
rect 2203 248 2205 250
rect 2199 247 2205 248
rect 2209 250 2215 251
rect 2209 248 2211 250
rect 2213 248 2215 250
rect 2237 249 2241 254
rect 2294 286 2307 287
rect 2294 284 2296 286
rect 2298 284 2307 286
rect 2294 283 2307 284
rect 2303 279 2319 283
rect 2291 275 2295 277
rect 1996 245 2021 246
rect 2105 245 2130 246
rect 2135 245 2139 247
rect 1987 243 1988 245
rect 1990 243 1991 245
rect 2135 243 2136 245
rect 2138 243 2139 245
rect 1987 240 1991 243
rect 2043 242 2049 243
rect 2043 240 2045 242
rect 2047 240 2049 242
rect 2077 242 2083 243
rect 2077 240 2079 242
rect 2081 240 2083 242
rect 2135 240 2139 243
rect 2155 243 2161 244
rect 2155 241 2157 243
rect 2159 241 2161 243
rect 2155 240 2161 241
rect 2174 243 2180 244
rect 2174 241 2176 243
rect 2178 241 2180 243
rect 2174 240 2180 241
rect 2209 240 2215 248
rect 2226 248 2241 249
rect 2226 246 2228 248
rect 2230 246 2241 248
rect 2226 245 2241 246
rect 2244 248 2248 250
rect 2244 246 2245 248
rect 2247 246 2248 248
rect 2267 274 2292 275
rect 2267 272 2269 274
rect 2271 273 2292 274
rect 2294 273 2295 275
rect 2271 272 2295 273
rect 2267 271 2295 272
rect 2267 251 2271 271
rect 2291 261 2295 271
rect 2311 266 2312 272
rect 2315 262 2319 279
rect 2291 259 2302 261
rect 2291 257 2299 259
rect 2301 257 2302 259
rect 2315 260 2320 262
rect 2315 258 2317 260
rect 2319 258 2320 260
rect 2291 255 2302 257
rect 2305 256 2320 258
rect 2305 254 2319 256
rect 2267 250 2273 251
rect 2267 248 2269 250
rect 2271 248 2273 250
rect 2267 247 2273 248
rect 2277 250 2283 251
rect 2277 248 2279 250
rect 2281 248 2283 250
rect 2305 249 2309 254
rect 2244 240 2248 246
rect 2277 240 2283 248
rect 2294 248 2309 249
rect 2294 246 2296 248
rect 2298 246 2309 248
rect 2294 245 2309 246
rect 2312 248 2316 250
rect 2312 246 2313 248
rect 2315 246 2316 248
rect 2312 240 2316 246
rect 99 221 103 224
rect 155 222 157 224
rect 159 222 161 224
rect 155 221 161 222
rect 189 222 191 224
rect 193 222 195 224
rect 189 221 195 222
rect 247 221 251 224
rect 99 219 100 221
rect 102 219 103 221
rect 247 219 248 221
rect 250 219 251 221
rect 267 223 273 224
rect 267 221 269 223
rect 271 221 273 223
rect 267 220 273 221
rect 286 223 292 224
rect 286 221 288 223
rect 290 221 292 223
rect 286 220 292 221
rect 366 221 370 224
rect 422 222 424 224
rect 426 222 428 224
rect 422 221 428 222
rect 456 222 458 224
rect 460 222 462 224
rect 456 221 462 222
rect 514 221 518 224
rect 366 219 367 221
rect 369 219 370 221
rect 514 219 515 221
rect 517 219 518 221
rect 534 223 540 224
rect 534 221 536 223
rect 538 221 540 223
rect 534 220 540 221
rect 553 223 559 224
rect 553 221 555 223
rect 557 221 559 223
rect 553 220 559 221
rect 633 221 637 224
rect 689 222 691 224
rect 693 222 695 224
rect 689 221 695 222
rect 723 222 725 224
rect 727 222 729 224
rect 723 221 729 222
rect 781 221 785 224
rect 633 219 634 221
rect 636 219 637 221
rect 781 219 782 221
rect 784 219 785 221
rect 801 223 807 224
rect 801 221 803 223
rect 805 221 807 223
rect 801 220 807 221
rect 820 223 826 224
rect 820 221 822 223
rect 824 221 826 223
rect 820 220 826 221
rect 900 221 904 224
rect 956 222 958 224
rect 960 222 962 224
rect 956 221 962 222
rect 990 222 992 224
rect 994 222 996 224
rect 990 221 996 222
rect 1048 221 1052 224
rect 900 219 901 221
rect 903 219 904 221
rect 1048 219 1049 221
rect 1051 219 1052 221
rect 1068 223 1074 224
rect 1068 221 1070 223
rect 1072 221 1074 223
rect 1068 220 1074 221
rect 1087 223 1093 224
rect 1087 221 1089 223
rect 1091 221 1093 223
rect 1087 220 1093 221
rect 1167 221 1171 224
rect 1223 222 1225 224
rect 1227 222 1229 224
rect 1223 221 1229 222
rect 1257 222 1259 224
rect 1261 222 1263 224
rect 1257 221 1263 222
rect 1315 221 1319 224
rect 1167 219 1168 221
rect 1170 219 1171 221
rect 1315 219 1316 221
rect 1318 219 1319 221
rect 1335 223 1341 224
rect 1335 221 1337 223
rect 1339 221 1341 223
rect 1335 220 1341 221
rect 1354 223 1360 224
rect 1354 221 1356 223
rect 1358 221 1360 223
rect 1354 220 1360 221
rect 1434 221 1438 224
rect 1490 222 1492 224
rect 1494 222 1496 224
rect 1490 221 1496 222
rect 1524 222 1526 224
rect 1528 222 1530 224
rect 1524 221 1530 222
rect 1582 221 1586 224
rect 1434 219 1435 221
rect 1437 219 1438 221
rect 1582 219 1583 221
rect 1585 219 1586 221
rect 1602 223 1608 224
rect 1602 221 1604 223
rect 1606 221 1608 223
rect 1602 220 1608 221
rect 1621 223 1627 224
rect 1621 221 1623 223
rect 1625 221 1627 223
rect 1621 220 1627 221
rect 1701 221 1705 224
rect 1757 222 1759 224
rect 1761 222 1763 224
rect 1757 221 1763 222
rect 1791 222 1793 224
rect 1795 222 1797 224
rect 1791 221 1797 222
rect 1849 221 1853 224
rect 1701 219 1702 221
rect 1704 219 1705 221
rect 1849 219 1850 221
rect 1852 219 1853 221
rect 1869 223 1875 224
rect 1869 221 1871 223
rect 1873 221 1875 223
rect 1869 220 1875 221
rect 1888 223 1894 224
rect 1888 221 1890 223
rect 1892 221 1894 223
rect 1888 220 1894 221
rect 8 217 28 218
rect 8 215 10 217
rect 12 215 28 217
rect 8 214 28 215
rect 24 210 28 214
rect 48 217 68 218
rect 48 215 50 217
rect 52 215 68 217
rect 48 214 68 215
rect 39 211 40 213
rect 24 206 36 210
rect 32 201 36 206
rect 32 199 33 201
rect 35 199 36 201
rect 32 187 36 199
rect 64 210 68 214
rect 79 211 80 213
rect 64 206 76 210
rect 72 201 76 206
rect 72 199 73 201
rect 75 199 76 201
rect 19 184 36 187
rect 19 182 20 184
rect 22 183 36 184
rect 22 182 23 183
rect 8 177 14 178
rect 8 175 10 177
rect 12 175 14 177
rect 8 168 14 175
rect 19 177 23 182
rect 72 187 76 199
rect 59 184 76 187
rect 59 182 60 184
rect 62 183 76 184
rect 62 182 63 183
rect 19 175 20 177
rect 22 175 23 177
rect 19 173 23 175
rect 28 179 34 180
rect 28 177 30 179
rect 32 177 34 179
rect 28 168 34 177
rect 48 177 54 178
rect 48 175 50 177
rect 52 175 54 177
rect 48 168 54 175
rect 59 177 63 182
rect 99 217 103 219
rect 108 218 133 219
rect 217 218 242 219
rect 108 216 110 218
rect 112 217 133 218
rect 112 216 130 217
rect 108 215 130 216
rect 132 215 133 217
rect 109 210 124 211
rect 109 209 120 210
rect 95 208 120 209
rect 122 208 124 210
rect 95 206 97 208
rect 99 207 124 208
rect 129 210 133 215
rect 138 217 148 218
rect 138 215 140 217
rect 142 215 148 217
rect 138 214 148 215
rect 129 208 130 210
rect 132 208 133 210
rect 99 206 113 207
rect 129 206 133 208
rect 95 205 113 206
rect 102 198 106 200
rect 102 196 103 198
rect 105 196 106 198
rect 102 186 106 196
rect 109 194 113 205
rect 144 210 148 214
rect 144 206 164 210
rect 160 203 164 206
rect 152 201 156 203
rect 152 199 153 201
rect 155 199 156 201
rect 152 194 156 199
rect 160 201 166 203
rect 160 199 163 201
rect 165 199 166 201
rect 160 197 166 199
rect 109 190 116 194
rect 112 189 116 190
rect 112 187 113 189
rect 115 187 116 189
rect 102 182 108 186
rect 112 185 116 187
rect 160 186 164 197
rect 124 185 164 186
rect 124 183 148 185
rect 150 183 164 185
rect 124 182 164 183
rect 59 175 60 177
rect 62 175 63 177
rect 59 173 63 175
rect 68 179 74 180
rect 68 177 70 179
rect 72 177 74 179
rect 104 178 128 182
rect 147 178 151 182
rect 202 217 212 218
rect 202 215 208 217
rect 210 215 212 217
rect 202 214 212 215
rect 217 217 238 218
rect 217 215 218 217
rect 220 216 238 217
rect 240 216 242 218
rect 247 217 251 219
rect 220 215 242 216
rect 202 210 206 214
rect 186 206 206 210
rect 186 203 190 206
rect 184 201 190 203
rect 184 199 185 201
rect 187 199 190 201
rect 184 197 190 199
rect 186 186 190 197
rect 194 201 198 203
rect 217 210 221 215
rect 315 217 335 218
rect 315 215 317 217
rect 319 215 335 217
rect 315 214 335 215
rect 217 208 218 210
rect 220 208 221 210
rect 217 206 221 208
rect 226 210 241 211
rect 226 208 228 210
rect 230 209 241 210
rect 230 208 255 209
rect 226 207 251 208
rect 237 206 251 207
rect 253 206 255 208
rect 237 205 255 206
rect 194 199 195 201
rect 197 199 198 201
rect 194 194 198 199
rect 237 194 241 205
rect 234 190 241 194
rect 244 198 248 200
rect 244 196 245 198
rect 247 196 248 198
rect 234 189 238 190
rect 234 187 235 189
rect 237 187 238 189
rect 186 185 226 186
rect 234 185 238 187
rect 244 186 248 196
rect 277 210 295 211
rect 277 208 279 210
rect 281 208 295 210
rect 277 207 295 208
rect 291 201 295 207
rect 291 199 292 201
rect 294 199 295 201
rect 270 194 276 195
rect 186 183 200 185
rect 202 183 226 185
rect 186 182 226 183
rect 242 182 248 186
rect 199 178 203 182
rect 222 178 246 182
rect 291 186 295 199
rect 280 182 295 186
rect 280 178 284 182
rect 298 178 299 189
rect 331 210 335 214
rect 346 211 347 213
rect 331 206 343 210
rect 339 201 343 206
rect 339 199 340 201
rect 342 199 343 201
rect 339 187 343 199
rect 326 184 343 187
rect 326 182 327 184
rect 329 183 343 184
rect 329 182 330 183
rect 68 168 74 177
rect 134 177 140 178
rect 134 175 136 177
rect 138 175 140 177
rect 99 170 105 171
rect 99 168 101 170
rect 103 168 105 170
rect 134 170 140 175
rect 147 176 148 178
rect 150 176 151 178
rect 147 174 151 176
rect 156 177 162 178
rect 156 175 158 177
rect 160 175 162 177
rect 134 168 136 170
rect 138 168 140 170
rect 156 170 162 175
rect 156 168 158 170
rect 160 168 162 170
rect 188 177 194 178
rect 188 175 190 177
rect 192 175 194 177
rect 188 170 194 175
rect 199 176 200 178
rect 202 176 203 178
rect 199 174 203 176
rect 210 177 216 178
rect 210 175 212 177
rect 214 175 216 177
rect 188 168 190 170
rect 192 168 194 170
rect 210 170 216 175
rect 267 177 284 178
rect 267 175 269 177
rect 271 175 284 177
rect 267 174 284 175
rect 315 177 321 178
rect 315 175 317 177
rect 319 175 321 177
rect 210 168 212 170
rect 214 168 216 170
rect 245 170 251 171
rect 245 168 247 170
rect 249 168 251 170
rect 286 170 292 171
rect 286 168 288 170
rect 290 168 292 170
rect 315 168 321 175
rect 326 177 330 182
rect 366 217 370 219
rect 375 218 400 219
rect 484 218 509 219
rect 375 216 377 218
rect 379 217 400 218
rect 379 216 397 217
rect 375 215 397 216
rect 399 215 400 217
rect 376 210 391 211
rect 376 209 387 210
rect 362 208 387 209
rect 389 208 391 210
rect 362 206 364 208
rect 366 207 391 208
rect 396 210 400 215
rect 405 217 415 218
rect 405 215 407 217
rect 409 215 415 217
rect 405 214 415 215
rect 396 208 397 210
rect 399 208 400 210
rect 366 206 380 207
rect 396 206 400 208
rect 362 205 380 206
rect 369 198 373 200
rect 369 196 370 198
rect 372 196 373 198
rect 369 186 373 196
rect 376 194 380 205
rect 411 210 415 214
rect 411 206 431 210
rect 427 203 431 206
rect 419 201 423 203
rect 419 199 420 201
rect 422 199 423 201
rect 419 194 423 199
rect 427 201 433 203
rect 427 199 430 201
rect 432 199 433 201
rect 427 197 433 199
rect 376 190 383 194
rect 379 189 383 190
rect 379 187 380 189
rect 382 187 383 189
rect 369 182 375 186
rect 379 185 383 187
rect 427 186 431 197
rect 391 185 431 186
rect 391 183 415 185
rect 417 183 431 185
rect 391 182 431 183
rect 326 175 327 177
rect 329 175 330 177
rect 326 173 330 175
rect 335 179 341 180
rect 335 177 337 179
rect 339 177 341 179
rect 371 178 395 182
rect 414 178 418 182
rect 469 217 479 218
rect 469 215 475 217
rect 477 215 479 217
rect 469 214 479 215
rect 484 217 505 218
rect 484 215 485 217
rect 487 216 505 217
rect 507 216 509 218
rect 514 217 518 219
rect 487 215 509 216
rect 469 210 473 214
rect 453 206 473 210
rect 453 203 457 206
rect 451 201 457 203
rect 451 199 452 201
rect 454 199 457 201
rect 451 197 457 199
rect 453 186 457 197
rect 461 201 465 203
rect 484 210 488 215
rect 582 217 602 218
rect 582 215 584 217
rect 586 215 602 217
rect 582 214 602 215
rect 484 208 485 210
rect 487 208 488 210
rect 484 206 488 208
rect 493 210 508 211
rect 493 208 495 210
rect 497 209 508 210
rect 497 208 522 209
rect 493 207 518 208
rect 504 206 518 207
rect 520 206 522 208
rect 504 205 522 206
rect 461 199 462 201
rect 464 199 465 201
rect 461 194 465 199
rect 504 194 508 205
rect 501 190 508 194
rect 511 198 515 200
rect 511 196 512 198
rect 514 196 515 198
rect 501 189 505 190
rect 501 187 502 189
rect 504 187 505 189
rect 453 185 493 186
rect 501 185 505 187
rect 511 186 515 196
rect 544 210 562 211
rect 544 208 546 210
rect 548 208 562 210
rect 544 207 562 208
rect 558 201 562 207
rect 558 199 559 201
rect 561 199 562 201
rect 537 194 543 195
rect 453 183 467 185
rect 469 183 493 185
rect 453 182 493 183
rect 509 182 515 186
rect 466 178 470 182
rect 489 178 513 182
rect 558 186 562 199
rect 547 182 562 186
rect 547 178 551 182
rect 565 178 566 189
rect 598 210 602 214
rect 613 211 614 213
rect 598 206 610 210
rect 606 201 610 206
rect 606 199 607 201
rect 609 199 610 201
rect 606 187 610 199
rect 593 184 610 187
rect 593 182 594 184
rect 596 183 610 184
rect 596 182 597 183
rect 335 168 341 177
rect 401 177 407 178
rect 401 175 403 177
rect 405 175 407 177
rect 366 170 372 171
rect 366 168 368 170
rect 370 168 372 170
rect 401 170 407 175
rect 414 176 415 178
rect 417 176 418 178
rect 414 174 418 176
rect 423 177 429 178
rect 423 175 425 177
rect 427 175 429 177
rect 401 168 403 170
rect 405 168 407 170
rect 423 170 429 175
rect 423 168 425 170
rect 427 168 429 170
rect 455 177 461 178
rect 455 175 457 177
rect 459 175 461 177
rect 455 170 461 175
rect 466 176 467 178
rect 469 176 470 178
rect 466 174 470 176
rect 477 177 483 178
rect 477 175 479 177
rect 481 175 483 177
rect 455 168 457 170
rect 459 168 461 170
rect 477 170 483 175
rect 534 177 551 178
rect 534 175 536 177
rect 538 175 551 177
rect 534 174 551 175
rect 582 177 588 178
rect 582 175 584 177
rect 586 175 588 177
rect 477 168 479 170
rect 481 168 483 170
rect 512 170 518 171
rect 512 168 514 170
rect 516 168 518 170
rect 553 170 559 171
rect 553 168 555 170
rect 557 168 559 170
rect 582 168 588 175
rect 593 177 597 182
rect 633 217 637 219
rect 642 218 667 219
rect 751 218 776 219
rect 642 216 644 218
rect 646 217 667 218
rect 646 216 664 217
rect 642 215 664 216
rect 666 215 667 217
rect 643 210 658 211
rect 643 209 654 210
rect 629 208 654 209
rect 656 208 658 210
rect 629 206 631 208
rect 633 207 658 208
rect 663 210 667 215
rect 672 217 682 218
rect 672 215 674 217
rect 676 215 682 217
rect 672 214 682 215
rect 663 208 664 210
rect 666 208 667 210
rect 633 206 647 207
rect 663 206 667 208
rect 629 205 647 206
rect 636 198 640 200
rect 636 196 637 198
rect 639 196 640 198
rect 636 186 640 196
rect 643 194 647 205
rect 678 210 682 214
rect 678 206 698 210
rect 694 203 698 206
rect 686 201 690 203
rect 686 199 687 201
rect 689 199 690 201
rect 686 194 690 199
rect 694 201 700 203
rect 694 199 697 201
rect 699 199 700 201
rect 694 197 700 199
rect 643 190 650 194
rect 646 189 650 190
rect 646 187 647 189
rect 649 187 650 189
rect 636 182 642 186
rect 646 185 650 187
rect 694 186 698 197
rect 658 185 698 186
rect 658 183 682 185
rect 684 183 698 185
rect 658 182 698 183
rect 593 175 594 177
rect 596 175 597 177
rect 593 173 597 175
rect 602 179 608 180
rect 602 177 604 179
rect 606 177 608 179
rect 638 178 662 182
rect 681 178 685 182
rect 736 217 746 218
rect 736 215 742 217
rect 744 215 746 217
rect 736 214 746 215
rect 751 217 772 218
rect 751 215 752 217
rect 754 216 772 217
rect 774 216 776 218
rect 781 217 785 219
rect 754 215 776 216
rect 736 210 740 214
rect 720 206 740 210
rect 720 203 724 206
rect 718 201 724 203
rect 718 199 719 201
rect 721 199 724 201
rect 718 197 724 199
rect 720 186 724 197
rect 728 201 732 203
rect 751 210 755 215
rect 849 217 869 218
rect 849 215 851 217
rect 853 215 869 217
rect 849 214 869 215
rect 751 208 752 210
rect 754 208 755 210
rect 751 206 755 208
rect 760 210 775 211
rect 760 208 762 210
rect 764 209 775 210
rect 764 208 789 209
rect 760 207 785 208
rect 771 206 785 207
rect 787 206 789 208
rect 771 205 789 206
rect 728 199 729 201
rect 731 199 732 201
rect 728 194 732 199
rect 771 194 775 205
rect 768 190 775 194
rect 778 198 782 200
rect 778 196 779 198
rect 781 196 782 198
rect 768 189 772 190
rect 768 187 769 189
rect 771 187 772 189
rect 720 185 760 186
rect 768 185 772 187
rect 778 186 782 196
rect 811 210 829 211
rect 811 208 813 210
rect 815 208 829 210
rect 811 207 829 208
rect 825 201 829 207
rect 825 199 826 201
rect 828 199 829 201
rect 804 194 810 195
rect 720 183 734 185
rect 736 183 760 185
rect 720 182 760 183
rect 776 182 782 186
rect 733 178 737 182
rect 756 178 780 182
rect 825 186 829 199
rect 814 182 829 186
rect 814 178 818 182
rect 832 178 833 189
rect 865 210 869 214
rect 880 211 881 213
rect 865 206 877 210
rect 873 201 877 206
rect 873 199 874 201
rect 876 199 877 201
rect 873 187 877 199
rect 860 184 877 187
rect 860 182 861 184
rect 863 183 877 184
rect 863 182 864 183
rect 602 168 608 177
rect 668 177 674 178
rect 668 175 670 177
rect 672 175 674 177
rect 633 170 639 171
rect 633 168 635 170
rect 637 168 639 170
rect 668 170 674 175
rect 681 176 682 178
rect 684 176 685 178
rect 681 174 685 176
rect 690 177 696 178
rect 690 175 692 177
rect 694 175 696 177
rect 668 168 670 170
rect 672 168 674 170
rect 690 170 696 175
rect 690 168 692 170
rect 694 168 696 170
rect 722 177 728 178
rect 722 175 724 177
rect 726 175 728 177
rect 722 170 728 175
rect 733 176 734 178
rect 736 176 737 178
rect 733 174 737 176
rect 744 177 750 178
rect 744 175 746 177
rect 748 175 750 177
rect 722 168 724 170
rect 726 168 728 170
rect 744 170 750 175
rect 801 177 818 178
rect 801 175 803 177
rect 805 175 818 177
rect 801 174 818 175
rect 849 177 855 178
rect 849 175 851 177
rect 853 175 855 177
rect 744 168 746 170
rect 748 168 750 170
rect 779 170 785 171
rect 779 168 781 170
rect 783 168 785 170
rect 820 170 826 171
rect 820 168 822 170
rect 824 168 826 170
rect 849 168 855 175
rect 860 177 864 182
rect 900 217 904 219
rect 909 218 934 219
rect 1018 218 1043 219
rect 909 216 911 218
rect 913 217 934 218
rect 913 216 931 217
rect 909 215 931 216
rect 933 215 934 217
rect 910 210 925 211
rect 910 209 921 210
rect 896 208 921 209
rect 923 208 925 210
rect 896 206 898 208
rect 900 207 925 208
rect 930 210 934 215
rect 939 217 949 218
rect 939 215 941 217
rect 943 215 949 217
rect 939 214 949 215
rect 930 208 931 210
rect 933 208 934 210
rect 900 206 914 207
rect 930 206 934 208
rect 896 205 914 206
rect 903 198 907 200
rect 903 196 904 198
rect 906 196 907 198
rect 903 186 907 196
rect 910 194 914 205
rect 945 210 949 214
rect 945 206 965 210
rect 961 203 965 206
rect 953 201 957 203
rect 953 199 954 201
rect 956 199 957 201
rect 953 194 957 199
rect 961 201 967 203
rect 961 199 964 201
rect 966 199 967 201
rect 961 197 967 199
rect 910 190 917 194
rect 913 189 917 190
rect 913 187 914 189
rect 916 187 917 189
rect 903 182 909 186
rect 913 185 917 187
rect 961 186 965 197
rect 925 185 965 186
rect 925 183 949 185
rect 951 183 965 185
rect 925 182 965 183
rect 860 175 861 177
rect 863 175 864 177
rect 860 173 864 175
rect 869 179 875 180
rect 869 177 871 179
rect 873 177 875 179
rect 905 178 929 182
rect 948 178 952 182
rect 1003 217 1013 218
rect 1003 215 1009 217
rect 1011 215 1013 217
rect 1003 214 1013 215
rect 1018 217 1039 218
rect 1018 215 1019 217
rect 1021 216 1039 217
rect 1041 216 1043 218
rect 1048 217 1052 219
rect 1021 215 1043 216
rect 1003 210 1007 214
rect 987 206 1007 210
rect 987 203 991 206
rect 985 201 991 203
rect 985 199 986 201
rect 988 199 991 201
rect 985 197 991 199
rect 987 186 991 197
rect 995 201 999 203
rect 1018 210 1022 215
rect 1116 217 1136 218
rect 1116 215 1118 217
rect 1120 215 1136 217
rect 1116 214 1136 215
rect 1018 208 1019 210
rect 1021 208 1022 210
rect 1018 206 1022 208
rect 1027 210 1042 211
rect 1027 208 1029 210
rect 1031 209 1042 210
rect 1031 208 1056 209
rect 1027 207 1052 208
rect 1038 206 1052 207
rect 1054 206 1056 208
rect 1038 205 1056 206
rect 995 199 996 201
rect 998 199 999 201
rect 995 194 999 199
rect 1038 194 1042 205
rect 1035 190 1042 194
rect 1045 198 1049 200
rect 1045 196 1046 198
rect 1048 196 1049 198
rect 1035 189 1039 190
rect 1035 187 1036 189
rect 1038 187 1039 189
rect 987 185 1027 186
rect 1035 185 1039 187
rect 1045 186 1049 196
rect 1078 210 1096 211
rect 1078 208 1080 210
rect 1082 208 1096 210
rect 1078 207 1096 208
rect 1092 201 1096 207
rect 1092 199 1093 201
rect 1095 199 1096 201
rect 1071 194 1077 195
rect 987 183 1001 185
rect 1003 183 1027 185
rect 987 182 1027 183
rect 1043 182 1049 186
rect 1000 178 1004 182
rect 1023 178 1047 182
rect 1092 186 1096 199
rect 1081 182 1096 186
rect 1081 178 1085 182
rect 1099 178 1100 189
rect 1132 210 1136 214
rect 1147 211 1148 213
rect 1132 206 1144 210
rect 1140 201 1144 206
rect 1140 199 1141 201
rect 1143 199 1144 201
rect 1140 187 1144 199
rect 1127 184 1144 187
rect 1127 182 1128 184
rect 1130 183 1144 184
rect 1130 182 1131 183
rect 869 168 875 177
rect 935 177 941 178
rect 935 175 937 177
rect 939 175 941 177
rect 900 170 906 171
rect 900 168 902 170
rect 904 168 906 170
rect 935 170 941 175
rect 948 176 949 178
rect 951 176 952 178
rect 948 174 952 176
rect 957 177 963 178
rect 957 175 959 177
rect 961 175 963 177
rect 935 168 937 170
rect 939 168 941 170
rect 957 170 963 175
rect 957 168 959 170
rect 961 168 963 170
rect 989 177 995 178
rect 989 175 991 177
rect 993 175 995 177
rect 989 170 995 175
rect 1000 176 1001 178
rect 1003 176 1004 178
rect 1000 174 1004 176
rect 1011 177 1017 178
rect 1011 175 1013 177
rect 1015 175 1017 177
rect 989 168 991 170
rect 993 168 995 170
rect 1011 170 1017 175
rect 1068 177 1085 178
rect 1068 175 1070 177
rect 1072 175 1085 177
rect 1068 174 1085 175
rect 1116 177 1122 178
rect 1116 175 1118 177
rect 1120 175 1122 177
rect 1011 168 1013 170
rect 1015 168 1017 170
rect 1046 170 1052 171
rect 1046 168 1048 170
rect 1050 168 1052 170
rect 1087 170 1093 171
rect 1087 168 1089 170
rect 1091 168 1093 170
rect 1116 168 1122 175
rect 1127 177 1131 182
rect 1167 217 1171 219
rect 1176 218 1201 219
rect 1285 218 1310 219
rect 1176 216 1178 218
rect 1180 217 1201 218
rect 1180 216 1198 217
rect 1176 215 1198 216
rect 1200 215 1201 217
rect 1177 210 1192 211
rect 1177 209 1188 210
rect 1163 208 1188 209
rect 1190 208 1192 210
rect 1163 206 1165 208
rect 1167 207 1192 208
rect 1197 210 1201 215
rect 1206 217 1216 218
rect 1206 215 1208 217
rect 1210 215 1216 217
rect 1206 214 1216 215
rect 1197 208 1198 210
rect 1200 208 1201 210
rect 1167 206 1181 207
rect 1197 206 1201 208
rect 1163 205 1181 206
rect 1170 198 1174 200
rect 1170 196 1171 198
rect 1173 196 1174 198
rect 1170 186 1174 196
rect 1177 194 1181 205
rect 1212 210 1216 214
rect 1212 206 1232 210
rect 1228 203 1232 206
rect 1220 201 1224 203
rect 1220 199 1221 201
rect 1223 199 1224 201
rect 1220 194 1224 199
rect 1228 201 1234 203
rect 1228 199 1231 201
rect 1233 199 1234 201
rect 1228 197 1234 199
rect 1177 190 1184 194
rect 1180 189 1184 190
rect 1180 187 1181 189
rect 1183 187 1184 189
rect 1170 182 1176 186
rect 1180 185 1184 187
rect 1228 186 1232 197
rect 1192 185 1232 186
rect 1192 183 1216 185
rect 1218 183 1232 185
rect 1192 182 1232 183
rect 1127 175 1128 177
rect 1130 175 1131 177
rect 1127 173 1131 175
rect 1136 179 1142 180
rect 1136 177 1138 179
rect 1140 177 1142 179
rect 1172 178 1196 182
rect 1215 178 1219 182
rect 1270 217 1280 218
rect 1270 215 1276 217
rect 1278 215 1280 217
rect 1270 214 1280 215
rect 1285 217 1306 218
rect 1285 215 1286 217
rect 1288 216 1306 217
rect 1308 216 1310 218
rect 1315 217 1319 219
rect 1288 215 1310 216
rect 1270 210 1274 214
rect 1254 206 1274 210
rect 1254 203 1258 206
rect 1252 201 1258 203
rect 1252 199 1253 201
rect 1255 199 1258 201
rect 1252 197 1258 199
rect 1254 186 1258 197
rect 1262 201 1266 203
rect 1285 210 1289 215
rect 1383 217 1403 218
rect 1383 215 1385 217
rect 1387 215 1403 217
rect 1383 214 1403 215
rect 1285 208 1286 210
rect 1288 208 1289 210
rect 1285 206 1289 208
rect 1294 210 1309 211
rect 1294 208 1296 210
rect 1298 209 1309 210
rect 1298 208 1323 209
rect 1294 207 1319 208
rect 1305 206 1319 207
rect 1321 206 1323 208
rect 1305 205 1323 206
rect 1262 199 1263 201
rect 1265 199 1266 201
rect 1262 194 1266 199
rect 1305 194 1309 205
rect 1302 190 1309 194
rect 1312 198 1316 200
rect 1312 196 1313 198
rect 1315 196 1316 198
rect 1302 189 1306 190
rect 1302 187 1303 189
rect 1305 187 1306 189
rect 1254 185 1294 186
rect 1302 185 1306 187
rect 1312 186 1316 196
rect 1345 210 1363 211
rect 1345 208 1347 210
rect 1349 208 1363 210
rect 1345 207 1363 208
rect 1359 201 1363 207
rect 1359 199 1360 201
rect 1362 199 1363 201
rect 1338 194 1344 195
rect 1254 183 1268 185
rect 1270 183 1294 185
rect 1254 182 1294 183
rect 1310 182 1316 186
rect 1267 178 1271 182
rect 1290 178 1314 182
rect 1359 186 1363 199
rect 1348 182 1363 186
rect 1348 178 1352 182
rect 1366 178 1367 189
rect 1399 210 1403 214
rect 1414 211 1415 213
rect 1399 206 1411 210
rect 1407 201 1411 206
rect 1407 199 1408 201
rect 1410 199 1411 201
rect 1407 187 1411 199
rect 1394 184 1411 187
rect 1394 182 1395 184
rect 1397 183 1411 184
rect 1397 182 1398 183
rect 1136 168 1142 177
rect 1202 177 1208 178
rect 1202 175 1204 177
rect 1206 175 1208 177
rect 1167 170 1173 171
rect 1167 168 1169 170
rect 1171 168 1173 170
rect 1202 170 1208 175
rect 1215 176 1216 178
rect 1218 176 1219 178
rect 1215 174 1219 176
rect 1224 177 1230 178
rect 1224 175 1226 177
rect 1228 175 1230 177
rect 1202 168 1204 170
rect 1206 168 1208 170
rect 1224 170 1230 175
rect 1224 168 1226 170
rect 1228 168 1230 170
rect 1256 177 1262 178
rect 1256 175 1258 177
rect 1260 175 1262 177
rect 1256 170 1262 175
rect 1267 176 1268 178
rect 1270 176 1271 178
rect 1267 174 1271 176
rect 1278 177 1284 178
rect 1278 175 1280 177
rect 1282 175 1284 177
rect 1256 168 1258 170
rect 1260 168 1262 170
rect 1278 170 1284 175
rect 1335 177 1352 178
rect 1335 175 1337 177
rect 1339 175 1352 177
rect 1335 174 1352 175
rect 1383 177 1389 178
rect 1383 175 1385 177
rect 1387 175 1389 177
rect 1278 168 1280 170
rect 1282 168 1284 170
rect 1313 170 1319 171
rect 1313 168 1315 170
rect 1317 168 1319 170
rect 1354 170 1360 171
rect 1354 168 1356 170
rect 1358 168 1360 170
rect 1383 168 1389 175
rect 1394 177 1398 182
rect 1434 217 1438 219
rect 1443 218 1468 219
rect 1552 218 1577 219
rect 1443 216 1445 218
rect 1447 217 1468 218
rect 1447 216 1465 217
rect 1443 215 1465 216
rect 1467 215 1468 217
rect 1444 210 1459 211
rect 1444 209 1455 210
rect 1430 208 1455 209
rect 1457 208 1459 210
rect 1430 206 1432 208
rect 1434 207 1459 208
rect 1464 210 1468 215
rect 1473 217 1483 218
rect 1473 215 1475 217
rect 1477 215 1483 217
rect 1473 214 1483 215
rect 1464 208 1465 210
rect 1467 208 1468 210
rect 1434 206 1448 207
rect 1464 206 1468 208
rect 1430 205 1448 206
rect 1437 198 1441 200
rect 1437 196 1438 198
rect 1440 196 1441 198
rect 1437 186 1441 196
rect 1444 194 1448 205
rect 1479 210 1483 214
rect 1479 206 1499 210
rect 1495 203 1499 206
rect 1487 201 1491 203
rect 1487 199 1488 201
rect 1490 199 1491 201
rect 1487 194 1491 199
rect 1495 201 1501 203
rect 1495 199 1498 201
rect 1500 199 1501 201
rect 1495 197 1501 199
rect 1444 190 1451 194
rect 1447 189 1451 190
rect 1447 187 1448 189
rect 1450 187 1451 189
rect 1437 182 1443 186
rect 1447 185 1451 187
rect 1495 186 1499 197
rect 1459 185 1499 186
rect 1459 183 1483 185
rect 1485 183 1499 185
rect 1459 182 1499 183
rect 1394 175 1395 177
rect 1397 175 1398 177
rect 1394 173 1398 175
rect 1403 179 1409 180
rect 1403 177 1405 179
rect 1407 177 1409 179
rect 1439 178 1463 182
rect 1482 178 1486 182
rect 1537 217 1547 218
rect 1537 215 1543 217
rect 1545 215 1547 217
rect 1537 214 1547 215
rect 1552 217 1573 218
rect 1552 215 1553 217
rect 1555 216 1573 217
rect 1575 216 1577 218
rect 1582 217 1586 219
rect 1555 215 1577 216
rect 1537 210 1541 214
rect 1521 206 1541 210
rect 1521 203 1525 206
rect 1519 201 1525 203
rect 1519 199 1520 201
rect 1522 199 1525 201
rect 1519 197 1525 199
rect 1521 186 1525 197
rect 1529 201 1533 203
rect 1552 210 1556 215
rect 1650 217 1670 218
rect 1650 215 1652 217
rect 1654 215 1670 217
rect 1650 214 1670 215
rect 1552 208 1553 210
rect 1555 208 1556 210
rect 1552 206 1556 208
rect 1561 210 1576 211
rect 1561 208 1563 210
rect 1565 209 1576 210
rect 1565 208 1590 209
rect 1561 207 1586 208
rect 1572 206 1586 207
rect 1588 206 1590 208
rect 1572 205 1590 206
rect 1529 199 1530 201
rect 1532 199 1533 201
rect 1529 194 1533 199
rect 1572 194 1576 205
rect 1569 190 1576 194
rect 1579 198 1583 200
rect 1579 196 1580 198
rect 1582 196 1583 198
rect 1569 189 1573 190
rect 1569 187 1570 189
rect 1572 187 1573 189
rect 1521 185 1561 186
rect 1569 185 1573 187
rect 1579 186 1583 196
rect 1612 210 1630 211
rect 1612 208 1614 210
rect 1616 208 1630 210
rect 1612 207 1630 208
rect 1626 201 1630 207
rect 1626 199 1627 201
rect 1629 199 1630 201
rect 1605 194 1611 195
rect 1521 183 1535 185
rect 1537 183 1561 185
rect 1521 182 1561 183
rect 1577 182 1583 186
rect 1534 178 1538 182
rect 1557 178 1581 182
rect 1626 186 1630 199
rect 1615 182 1630 186
rect 1615 178 1619 182
rect 1633 178 1634 189
rect 1666 210 1670 214
rect 1681 211 1682 213
rect 1666 206 1678 210
rect 1674 201 1678 206
rect 1674 199 1675 201
rect 1677 199 1678 201
rect 1674 187 1678 199
rect 1661 184 1678 187
rect 1661 182 1662 184
rect 1664 183 1678 184
rect 1664 182 1665 183
rect 1403 168 1409 177
rect 1469 177 1475 178
rect 1469 175 1471 177
rect 1473 175 1475 177
rect 1434 170 1440 171
rect 1434 168 1436 170
rect 1438 168 1440 170
rect 1469 170 1475 175
rect 1482 176 1483 178
rect 1485 176 1486 178
rect 1482 174 1486 176
rect 1491 177 1497 178
rect 1491 175 1493 177
rect 1495 175 1497 177
rect 1469 168 1471 170
rect 1473 168 1475 170
rect 1491 170 1497 175
rect 1491 168 1493 170
rect 1495 168 1497 170
rect 1523 177 1529 178
rect 1523 175 1525 177
rect 1527 175 1529 177
rect 1523 170 1529 175
rect 1534 176 1535 178
rect 1537 176 1538 178
rect 1534 174 1538 176
rect 1545 177 1551 178
rect 1545 175 1547 177
rect 1549 175 1551 177
rect 1523 168 1525 170
rect 1527 168 1529 170
rect 1545 170 1551 175
rect 1602 177 1619 178
rect 1602 175 1604 177
rect 1606 175 1619 177
rect 1602 174 1619 175
rect 1650 177 1656 178
rect 1650 175 1652 177
rect 1654 175 1656 177
rect 1545 168 1547 170
rect 1549 168 1551 170
rect 1580 170 1586 171
rect 1580 168 1582 170
rect 1584 168 1586 170
rect 1621 170 1627 171
rect 1621 168 1623 170
rect 1625 168 1627 170
rect 1650 168 1656 175
rect 1661 177 1665 182
rect 1701 217 1705 219
rect 1710 218 1735 219
rect 1819 218 1844 219
rect 1710 216 1712 218
rect 1714 217 1735 218
rect 1714 216 1732 217
rect 1710 215 1732 216
rect 1734 215 1735 217
rect 1711 210 1726 211
rect 1711 209 1722 210
rect 1697 208 1722 209
rect 1724 208 1726 210
rect 1697 206 1699 208
rect 1701 207 1726 208
rect 1731 210 1735 215
rect 1740 217 1750 218
rect 1740 215 1742 217
rect 1744 215 1750 217
rect 1740 214 1750 215
rect 1731 208 1732 210
rect 1734 208 1735 210
rect 1701 206 1715 207
rect 1731 206 1735 208
rect 1697 205 1715 206
rect 1704 198 1708 200
rect 1704 196 1705 198
rect 1707 196 1708 198
rect 1704 186 1708 196
rect 1711 194 1715 205
rect 1746 210 1750 214
rect 1746 206 1766 210
rect 1762 203 1766 206
rect 1754 201 1758 203
rect 1754 199 1755 201
rect 1757 199 1758 201
rect 1754 194 1758 199
rect 1762 201 1768 203
rect 1762 199 1765 201
rect 1767 199 1768 201
rect 1762 197 1768 199
rect 1711 190 1718 194
rect 1714 189 1718 190
rect 1714 187 1715 189
rect 1717 187 1718 189
rect 1704 182 1710 186
rect 1714 185 1718 187
rect 1762 186 1766 197
rect 1726 185 1766 186
rect 1726 183 1750 185
rect 1752 183 1766 185
rect 1726 182 1766 183
rect 1661 175 1662 177
rect 1664 175 1665 177
rect 1661 173 1665 175
rect 1670 179 1676 180
rect 1670 177 1672 179
rect 1674 177 1676 179
rect 1706 178 1730 182
rect 1749 178 1753 182
rect 1804 217 1814 218
rect 1804 215 1810 217
rect 1812 215 1814 217
rect 1804 214 1814 215
rect 1819 217 1840 218
rect 1819 215 1820 217
rect 1822 216 1840 217
rect 1842 216 1844 218
rect 1849 217 1853 219
rect 1822 215 1844 216
rect 1926 218 1932 224
rect 1987 221 1991 224
rect 2043 222 2045 224
rect 2047 222 2049 224
rect 2043 221 2049 222
rect 2077 222 2079 224
rect 2081 222 2083 224
rect 2077 221 2083 222
rect 2135 221 2139 224
rect 1987 219 1988 221
rect 1990 219 1991 221
rect 2135 219 2136 221
rect 2138 219 2139 221
rect 2155 223 2161 224
rect 2155 221 2157 223
rect 2159 221 2161 223
rect 2155 220 2161 221
rect 2174 223 2180 224
rect 2174 221 2176 223
rect 2178 221 2180 223
rect 2174 220 2180 221
rect 1926 216 1928 218
rect 1930 216 1932 218
rect 1926 215 1932 216
rect 1939 215 1943 217
rect 1804 210 1808 214
rect 1788 206 1808 210
rect 1788 203 1792 206
rect 1786 201 1792 203
rect 1786 199 1787 201
rect 1789 199 1792 201
rect 1786 197 1792 199
rect 1788 186 1792 197
rect 1796 201 1800 203
rect 1819 210 1823 215
rect 1939 213 1940 215
rect 1942 213 1943 215
rect 1819 208 1820 210
rect 1822 208 1823 210
rect 1819 206 1823 208
rect 1828 210 1843 211
rect 1828 208 1830 210
rect 1832 209 1843 210
rect 1832 208 1857 209
rect 1828 207 1853 208
rect 1839 206 1853 207
rect 1855 206 1857 208
rect 1839 205 1857 206
rect 1796 199 1797 201
rect 1799 199 1800 201
rect 1796 194 1800 199
rect 1839 194 1843 205
rect 1836 190 1843 194
rect 1846 198 1850 200
rect 1846 196 1847 198
rect 1849 196 1850 198
rect 1836 189 1840 190
rect 1836 187 1837 189
rect 1839 187 1840 189
rect 1788 185 1828 186
rect 1836 185 1840 187
rect 1846 186 1850 196
rect 1879 210 1897 211
rect 1879 208 1881 210
rect 1883 208 1897 210
rect 1879 207 1897 208
rect 1893 201 1897 207
rect 1893 199 1894 201
rect 1896 199 1897 201
rect 1872 194 1878 195
rect 1788 183 1802 185
rect 1804 183 1828 185
rect 1788 182 1828 183
rect 1844 182 1850 186
rect 1801 178 1805 182
rect 1824 178 1848 182
rect 1893 186 1897 199
rect 1882 182 1897 186
rect 1882 178 1886 182
rect 1900 178 1901 189
rect 1913 210 1917 212
rect 1913 208 1914 210
rect 1916 208 1917 210
rect 1913 202 1917 208
rect 1939 210 1943 213
rect 1939 206 1963 210
rect 1913 198 1924 202
rect 1670 168 1676 177
rect 1736 177 1742 178
rect 1736 175 1738 177
rect 1740 175 1742 177
rect 1701 170 1707 171
rect 1701 168 1703 170
rect 1705 168 1707 170
rect 1736 170 1742 175
rect 1749 176 1750 178
rect 1752 176 1753 178
rect 1749 174 1753 176
rect 1758 177 1764 178
rect 1758 175 1760 177
rect 1762 175 1764 177
rect 1736 168 1738 170
rect 1740 168 1742 170
rect 1758 170 1764 175
rect 1758 168 1760 170
rect 1762 168 1764 170
rect 1790 177 1796 178
rect 1790 175 1792 177
rect 1794 175 1796 177
rect 1790 170 1796 175
rect 1801 176 1802 178
rect 1804 176 1805 178
rect 1801 174 1805 176
rect 1812 177 1818 178
rect 1812 175 1814 177
rect 1816 175 1818 177
rect 1790 168 1792 170
rect 1794 168 1796 170
rect 1812 170 1818 175
rect 1869 177 1886 178
rect 1869 175 1871 177
rect 1873 175 1886 177
rect 1869 174 1886 175
rect 1920 192 1924 198
rect 1959 202 1963 206
rect 1939 201 1955 202
rect 1939 199 1951 201
rect 1953 199 1955 201
rect 1939 198 1955 199
rect 1959 200 1964 202
rect 1959 198 1961 200
rect 1963 198 1964 200
rect 1939 192 1943 198
rect 1959 196 1964 198
rect 1959 194 1963 196
rect 1920 191 1943 192
rect 1920 189 1922 191
rect 1924 189 1943 191
rect 1920 188 1943 189
rect 1931 177 1935 179
rect 1931 175 1932 177
rect 1934 175 1935 177
rect 1812 168 1814 170
rect 1816 168 1818 170
rect 1847 170 1853 171
rect 1847 168 1849 170
rect 1851 168 1853 170
rect 1888 170 1894 171
rect 1888 168 1890 170
rect 1892 168 1894 170
rect 1931 170 1935 175
rect 1939 177 1943 188
rect 1947 191 1963 194
rect 1947 189 1948 191
rect 1950 190 1963 191
rect 1950 189 1951 190
rect 1947 184 1951 189
rect 1947 182 1948 184
rect 1950 182 1951 184
rect 1947 180 1951 182
rect 1987 217 1991 219
rect 1996 218 2021 219
rect 2105 218 2130 219
rect 1996 216 1998 218
rect 2000 217 2021 218
rect 2000 216 2018 217
rect 1996 215 2018 216
rect 2020 215 2021 217
rect 1997 210 2012 211
rect 1997 209 2008 210
rect 1983 208 2008 209
rect 2010 208 2012 210
rect 1983 206 1985 208
rect 1987 207 2012 208
rect 2017 210 2021 215
rect 2026 217 2036 218
rect 2026 215 2028 217
rect 2030 215 2036 217
rect 2026 214 2036 215
rect 2017 208 2018 210
rect 2020 208 2021 210
rect 1987 206 2001 207
rect 2017 206 2021 208
rect 1983 205 2001 206
rect 1990 198 1994 200
rect 1990 196 1991 198
rect 1993 196 1994 198
rect 1990 186 1994 196
rect 1997 194 2001 205
rect 2032 210 2036 214
rect 2032 206 2052 210
rect 2048 203 2052 206
rect 2040 201 2044 203
rect 2040 199 2041 201
rect 2043 199 2044 201
rect 2040 194 2044 199
rect 2048 201 2054 203
rect 2048 199 2051 201
rect 2053 199 2054 201
rect 2048 197 2054 199
rect 1997 190 2004 194
rect 2000 189 2004 190
rect 2000 187 2001 189
rect 2003 187 2004 189
rect 1990 182 1996 186
rect 2000 185 2004 187
rect 2048 186 2052 197
rect 2012 185 2052 186
rect 2012 183 2036 185
rect 2038 183 2052 185
rect 2012 182 2052 183
rect 1992 178 2016 182
rect 2035 178 2039 182
rect 2090 217 2100 218
rect 2090 215 2096 217
rect 2098 215 2100 217
rect 2090 214 2100 215
rect 2105 217 2126 218
rect 2105 215 2106 217
rect 2108 216 2126 217
rect 2128 216 2130 218
rect 2135 217 2139 219
rect 2108 215 2130 216
rect 2199 216 2205 217
rect 2090 210 2094 214
rect 2074 206 2094 210
rect 2074 203 2078 206
rect 2072 201 2078 203
rect 2072 199 2073 201
rect 2075 199 2078 201
rect 2072 197 2078 199
rect 2074 186 2078 197
rect 2082 201 2086 203
rect 2105 210 2109 215
rect 2105 208 2106 210
rect 2108 208 2109 210
rect 2105 206 2109 208
rect 2114 210 2129 211
rect 2114 208 2116 210
rect 2118 209 2129 210
rect 2118 208 2143 209
rect 2114 207 2139 208
rect 2125 206 2139 207
rect 2141 206 2143 208
rect 2125 205 2143 206
rect 2082 199 2083 201
rect 2085 199 2086 201
rect 2082 194 2086 199
rect 2125 194 2129 205
rect 2122 190 2129 194
rect 2132 198 2136 200
rect 2132 196 2133 198
rect 2135 196 2136 198
rect 2122 189 2126 190
rect 2122 187 2123 189
rect 2125 187 2126 189
rect 2074 185 2114 186
rect 2122 185 2126 187
rect 2132 186 2136 196
rect 2199 214 2201 216
rect 2203 214 2205 216
rect 2199 213 2205 214
rect 2209 216 2215 224
rect 2209 214 2211 216
rect 2213 214 2215 216
rect 2226 218 2241 219
rect 2226 216 2228 218
rect 2230 216 2241 218
rect 2226 215 2241 216
rect 2209 213 2215 214
rect 2165 210 2183 211
rect 2165 208 2167 210
rect 2169 208 2183 210
rect 2165 207 2183 208
rect 2179 201 2183 207
rect 2179 199 2180 201
rect 2182 199 2183 201
rect 2158 194 2164 195
rect 2074 183 2088 185
rect 2090 183 2114 185
rect 2074 182 2114 183
rect 2130 182 2136 186
rect 2087 178 2091 182
rect 2110 178 2134 182
rect 2179 186 2183 199
rect 2168 182 2183 186
rect 2168 178 2172 182
rect 2186 178 2187 189
rect 2199 193 2203 213
rect 2237 210 2241 215
rect 2244 218 2248 224
rect 2244 216 2245 218
rect 2247 216 2248 218
rect 2244 214 2248 216
rect 2223 207 2234 209
rect 2223 205 2231 207
rect 2233 205 2234 207
rect 2237 208 2251 210
rect 2237 206 2252 208
rect 2223 203 2234 205
rect 2247 204 2249 206
rect 2251 204 2252 206
rect 2223 193 2227 203
rect 2247 202 2252 204
rect 2199 192 2227 193
rect 2199 190 2201 192
rect 2203 191 2227 192
rect 2203 190 2224 191
rect 2199 189 2224 190
rect 2226 189 2227 191
rect 2243 192 2244 198
rect 2223 187 2227 189
rect 2022 177 2028 178
rect 1939 176 1972 177
rect 1939 174 1968 176
rect 1970 174 1972 176
rect 1939 173 1972 174
rect 2022 175 2024 177
rect 2026 175 2028 177
rect 1931 168 1932 170
rect 1934 168 1935 170
rect 1987 170 1993 171
rect 1987 168 1989 170
rect 1991 168 1993 170
rect 2022 170 2028 175
rect 2035 176 2036 178
rect 2038 176 2039 178
rect 2035 174 2039 176
rect 2044 177 2050 178
rect 2044 175 2046 177
rect 2048 175 2050 177
rect 2022 168 2024 170
rect 2026 168 2028 170
rect 2044 170 2050 175
rect 2044 168 2046 170
rect 2048 168 2050 170
rect 2076 177 2082 178
rect 2076 175 2078 177
rect 2080 175 2082 177
rect 2076 170 2082 175
rect 2087 176 2088 178
rect 2090 176 2091 178
rect 2087 174 2091 176
rect 2098 177 2104 178
rect 2098 175 2100 177
rect 2102 175 2104 177
rect 2076 168 2078 170
rect 2080 168 2082 170
rect 2098 170 2104 175
rect 2155 177 2172 178
rect 2155 175 2157 177
rect 2159 175 2172 177
rect 2155 174 2172 175
rect 2247 185 2251 202
rect 2235 181 2251 185
rect 2226 180 2239 181
rect 2226 178 2228 180
rect 2230 178 2239 180
rect 2267 216 2273 217
rect 2267 214 2269 216
rect 2271 214 2273 216
rect 2267 213 2273 214
rect 2277 216 2283 224
rect 2277 214 2279 216
rect 2281 214 2283 216
rect 2294 218 2309 219
rect 2294 216 2296 218
rect 2298 216 2309 218
rect 2294 215 2309 216
rect 2277 213 2283 214
rect 2267 193 2271 213
rect 2305 210 2309 215
rect 2312 218 2316 224
rect 2312 216 2313 218
rect 2315 216 2316 218
rect 2312 214 2316 216
rect 2291 207 2302 209
rect 2291 205 2299 207
rect 2301 205 2302 207
rect 2305 208 2319 210
rect 2305 206 2320 208
rect 2291 203 2302 205
rect 2315 204 2317 206
rect 2319 204 2320 206
rect 2291 193 2295 203
rect 2315 202 2320 204
rect 2267 192 2295 193
rect 2267 190 2269 192
rect 2271 191 2295 192
rect 2271 190 2292 191
rect 2267 189 2292 190
rect 2294 189 2295 191
rect 2311 192 2312 198
rect 2291 187 2295 189
rect 2226 177 2239 178
rect 2315 185 2319 202
rect 2303 181 2319 185
rect 2294 180 2307 181
rect 2294 178 2296 180
rect 2298 178 2307 180
rect 2294 177 2307 178
rect 2098 168 2100 170
rect 2102 168 2104 170
rect 2133 170 2139 171
rect 2133 168 2135 170
rect 2137 168 2139 170
rect 2174 170 2180 171
rect 2174 168 2176 170
rect 2178 168 2180 170
rect 2210 170 2214 172
rect 2210 168 2211 170
rect 2213 168 2214 170
rect 2243 170 2249 171
rect 2243 168 2245 170
rect 2247 168 2249 170
rect 2278 170 2282 172
rect 2278 168 2279 170
rect 2281 168 2282 170
rect 2311 170 2317 171
rect 2311 168 2313 170
rect 2315 168 2317 170
rect 8 145 14 152
rect 8 143 10 145
rect 12 143 14 145
rect 8 142 14 143
rect 19 145 23 147
rect 19 143 20 145
rect 22 143 23 145
rect 19 138 23 143
rect 28 143 34 152
rect 48 145 54 152
rect 48 143 50 145
rect 52 143 54 145
rect 28 141 30 143
rect 32 141 34 143
rect 28 140 34 141
rect 48 142 54 143
rect 59 145 63 147
rect 59 143 60 145
rect 62 143 63 145
rect 19 136 20 138
rect 22 137 23 138
rect 22 136 36 137
rect 19 133 36 136
rect 32 121 36 133
rect 59 138 63 143
rect 68 143 74 152
rect 99 150 101 152
rect 103 150 105 152
rect 99 149 105 150
rect 134 150 136 152
rect 138 150 140 152
rect 68 141 70 143
rect 72 141 74 143
rect 134 145 140 150
rect 156 150 158 152
rect 160 150 162 152
rect 134 143 136 145
rect 138 143 140 145
rect 134 142 140 143
rect 147 144 151 146
rect 147 142 148 144
rect 150 142 151 144
rect 156 145 162 150
rect 156 143 158 145
rect 160 143 162 145
rect 156 142 162 143
rect 188 150 190 152
rect 192 150 194 152
rect 188 145 194 150
rect 210 150 212 152
rect 214 150 216 152
rect 188 143 190 145
rect 192 143 194 145
rect 188 142 194 143
rect 199 144 203 146
rect 199 142 200 144
rect 202 142 203 144
rect 210 145 216 150
rect 245 150 247 152
rect 249 150 251 152
rect 245 149 251 150
rect 286 150 288 152
rect 290 150 292 152
rect 286 149 292 150
rect 210 143 212 145
rect 214 143 216 145
rect 210 142 216 143
rect 267 145 284 146
rect 267 143 269 145
rect 271 143 284 145
rect 267 142 284 143
rect 315 145 321 152
rect 315 143 317 145
rect 319 143 321 145
rect 315 142 321 143
rect 326 145 330 147
rect 326 143 327 145
rect 329 143 330 145
rect 68 140 74 141
rect 59 136 60 138
rect 62 137 63 138
rect 62 136 76 137
rect 59 133 76 136
rect 32 119 33 121
rect 35 119 36 121
rect 32 114 36 119
rect 24 110 36 114
rect 24 106 28 110
rect 39 107 40 109
rect 72 121 76 133
rect 72 119 73 121
rect 75 119 76 121
rect 72 114 76 119
rect 64 110 76 114
rect 8 105 28 106
rect 8 103 10 105
rect 12 103 28 105
rect 8 102 28 103
rect 64 106 68 110
rect 79 107 80 109
rect 48 105 68 106
rect 48 103 50 105
rect 52 103 68 105
rect 48 102 68 103
rect 104 138 128 142
rect 147 138 151 142
rect 102 134 108 138
rect 124 137 164 138
rect 124 135 148 137
rect 150 135 164 137
rect 102 124 106 134
rect 112 133 116 135
rect 124 134 164 135
rect 112 131 113 133
rect 115 131 116 133
rect 112 130 116 131
rect 102 122 103 124
rect 105 122 106 124
rect 102 120 106 122
rect 109 126 116 130
rect 109 115 113 126
rect 152 121 156 126
rect 152 119 153 121
rect 155 119 156 121
rect 95 114 113 115
rect 95 112 97 114
rect 99 113 113 114
rect 99 112 124 113
rect 95 111 120 112
rect 109 110 120 111
rect 122 110 124 112
rect 109 109 124 110
rect 129 112 133 114
rect 129 110 130 112
rect 132 110 133 112
rect 129 105 133 110
rect 152 117 156 119
rect 160 123 164 134
rect 160 121 166 123
rect 160 119 163 121
rect 165 119 166 121
rect 160 117 166 119
rect 160 114 164 117
rect 144 110 164 114
rect 144 106 148 110
rect 108 104 130 105
rect 99 101 103 103
rect 108 102 110 104
rect 112 103 130 104
rect 132 103 133 105
rect 112 102 133 103
rect 138 105 148 106
rect 138 103 140 105
rect 142 103 148 105
rect 138 102 148 103
rect 199 138 203 142
rect 222 138 246 142
rect 186 137 226 138
rect 186 135 200 137
rect 202 135 226 137
rect 186 134 226 135
rect 186 123 190 134
rect 234 133 238 135
rect 242 134 248 138
rect 234 131 235 133
rect 237 131 238 133
rect 234 130 238 131
rect 234 126 241 130
rect 184 121 190 123
rect 184 119 185 121
rect 187 119 190 121
rect 184 117 190 119
rect 194 121 198 126
rect 194 119 195 121
rect 197 119 198 121
rect 194 117 198 119
rect 186 114 190 117
rect 186 110 206 114
rect 202 106 206 110
rect 237 115 241 126
rect 244 124 248 134
rect 244 122 245 124
rect 247 122 248 124
rect 244 120 248 122
rect 237 114 255 115
rect 217 112 221 114
rect 237 113 251 114
rect 217 110 218 112
rect 220 110 221 112
rect 202 105 212 106
rect 202 103 208 105
rect 210 103 212 105
rect 202 102 212 103
rect 217 105 221 110
rect 226 112 251 113
rect 253 112 255 114
rect 226 110 228 112
rect 230 111 255 112
rect 230 110 241 111
rect 226 109 241 110
rect 280 138 284 142
rect 280 134 295 138
rect 270 125 276 126
rect 291 121 295 134
rect 298 131 299 142
rect 291 119 292 121
rect 294 119 295 121
rect 291 113 295 119
rect 326 138 330 143
rect 335 143 341 152
rect 366 150 368 152
rect 370 150 372 152
rect 366 149 372 150
rect 401 150 403 152
rect 405 150 407 152
rect 335 141 337 143
rect 339 141 341 143
rect 401 145 407 150
rect 423 150 425 152
rect 427 150 429 152
rect 401 143 403 145
rect 405 143 407 145
rect 401 142 407 143
rect 414 144 418 146
rect 414 142 415 144
rect 417 142 418 144
rect 423 145 429 150
rect 423 143 425 145
rect 427 143 429 145
rect 423 142 429 143
rect 455 150 457 152
rect 459 150 461 152
rect 455 145 461 150
rect 477 150 479 152
rect 481 150 483 152
rect 455 143 457 145
rect 459 143 461 145
rect 455 142 461 143
rect 466 144 470 146
rect 466 142 467 144
rect 469 142 470 144
rect 477 145 483 150
rect 512 150 514 152
rect 516 150 518 152
rect 512 149 518 150
rect 553 150 555 152
rect 557 150 559 152
rect 553 149 559 150
rect 477 143 479 145
rect 481 143 483 145
rect 477 142 483 143
rect 534 145 551 146
rect 534 143 536 145
rect 538 143 551 145
rect 534 142 551 143
rect 582 145 588 152
rect 582 143 584 145
rect 586 143 588 145
rect 582 142 588 143
rect 593 145 597 147
rect 593 143 594 145
rect 596 143 597 145
rect 335 140 341 141
rect 326 136 327 138
rect 329 137 330 138
rect 329 136 343 137
rect 326 133 343 136
rect 277 112 295 113
rect 277 110 279 112
rect 281 110 295 112
rect 277 109 295 110
rect 339 121 343 133
rect 339 119 340 121
rect 342 119 343 121
rect 339 114 343 119
rect 331 110 343 114
rect 331 106 335 110
rect 346 107 347 109
rect 217 103 218 105
rect 220 104 242 105
rect 220 103 238 104
rect 217 102 238 103
rect 240 102 242 104
rect 108 101 133 102
rect 217 101 242 102
rect 247 101 251 103
rect 315 105 335 106
rect 315 103 317 105
rect 319 103 335 105
rect 315 102 335 103
rect 371 138 395 142
rect 414 138 418 142
rect 369 134 375 138
rect 391 137 431 138
rect 391 135 415 137
rect 417 135 431 137
rect 369 124 373 134
rect 379 133 383 135
rect 391 134 431 135
rect 379 131 380 133
rect 382 131 383 133
rect 379 130 383 131
rect 369 122 370 124
rect 372 122 373 124
rect 369 120 373 122
rect 376 126 383 130
rect 376 115 380 126
rect 419 121 423 126
rect 419 119 420 121
rect 422 119 423 121
rect 362 114 380 115
rect 362 112 364 114
rect 366 113 380 114
rect 366 112 391 113
rect 362 111 387 112
rect 376 110 387 111
rect 389 110 391 112
rect 376 109 391 110
rect 396 112 400 114
rect 396 110 397 112
rect 399 110 400 112
rect 396 105 400 110
rect 419 117 423 119
rect 427 123 431 134
rect 427 121 433 123
rect 427 119 430 121
rect 432 119 433 121
rect 427 117 433 119
rect 427 114 431 117
rect 411 110 431 114
rect 411 106 415 110
rect 375 104 397 105
rect 366 101 370 103
rect 375 102 377 104
rect 379 103 397 104
rect 399 103 400 105
rect 379 102 400 103
rect 405 105 415 106
rect 405 103 407 105
rect 409 103 415 105
rect 405 102 415 103
rect 466 138 470 142
rect 489 138 513 142
rect 453 137 493 138
rect 453 135 467 137
rect 469 135 493 137
rect 453 134 493 135
rect 453 123 457 134
rect 501 133 505 135
rect 509 134 515 138
rect 501 131 502 133
rect 504 131 505 133
rect 501 130 505 131
rect 501 126 508 130
rect 451 121 457 123
rect 451 119 452 121
rect 454 119 457 121
rect 451 117 457 119
rect 461 121 465 126
rect 461 119 462 121
rect 464 119 465 121
rect 461 117 465 119
rect 453 114 457 117
rect 453 110 473 114
rect 469 106 473 110
rect 504 115 508 126
rect 511 124 515 134
rect 511 122 512 124
rect 514 122 515 124
rect 511 120 515 122
rect 504 114 522 115
rect 484 112 488 114
rect 504 113 518 114
rect 484 110 485 112
rect 487 110 488 112
rect 469 105 479 106
rect 469 103 475 105
rect 477 103 479 105
rect 469 102 479 103
rect 484 105 488 110
rect 493 112 518 113
rect 520 112 522 114
rect 493 110 495 112
rect 497 111 522 112
rect 497 110 508 111
rect 493 109 508 110
rect 547 138 551 142
rect 547 134 562 138
rect 537 125 543 126
rect 558 121 562 134
rect 565 131 566 142
rect 558 119 559 121
rect 561 119 562 121
rect 558 113 562 119
rect 593 138 597 143
rect 602 143 608 152
rect 633 150 635 152
rect 637 150 639 152
rect 633 149 639 150
rect 668 150 670 152
rect 672 150 674 152
rect 602 141 604 143
rect 606 141 608 143
rect 668 145 674 150
rect 690 150 692 152
rect 694 150 696 152
rect 668 143 670 145
rect 672 143 674 145
rect 668 142 674 143
rect 681 144 685 146
rect 681 142 682 144
rect 684 142 685 144
rect 690 145 696 150
rect 690 143 692 145
rect 694 143 696 145
rect 690 142 696 143
rect 722 150 724 152
rect 726 150 728 152
rect 722 145 728 150
rect 744 150 746 152
rect 748 150 750 152
rect 722 143 724 145
rect 726 143 728 145
rect 722 142 728 143
rect 733 144 737 146
rect 733 142 734 144
rect 736 142 737 144
rect 744 145 750 150
rect 779 150 781 152
rect 783 150 785 152
rect 779 149 785 150
rect 820 150 822 152
rect 824 150 826 152
rect 820 149 826 150
rect 744 143 746 145
rect 748 143 750 145
rect 744 142 750 143
rect 801 145 818 146
rect 801 143 803 145
rect 805 143 818 145
rect 801 142 818 143
rect 849 145 855 152
rect 849 143 851 145
rect 853 143 855 145
rect 849 142 855 143
rect 860 145 864 147
rect 860 143 861 145
rect 863 143 864 145
rect 602 140 608 141
rect 593 136 594 138
rect 596 137 597 138
rect 596 136 610 137
rect 593 133 610 136
rect 544 112 562 113
rect 544 110 546 112
rect 548 110 562 112
rect 544 109 562 110
rect 606 121 610 133
rect 606 119 607 121
rect 609 119 610 121
rect 606 114 610 119
rect 598 110 610 114
rect 598 106 602 110
rect 613 107 614 109
rect 484 103 485 105
rect 487 104 509 105
rect 487 103 505 104
rect 484 102 505 103
rect 507 102 509 104
rect 375 101 400 102
rect 484 101 509 102
rect 514 101 518 103
rect 582 105 602 106
rect 582 103 584 105
rect 586 103 602 105
rect 582 102 602 103
rect 638 138 662 142
rect 681 138 685 142
rect 636 134 642 138
rect 658 137 698 138
rect 658 135 682 137
rect 684 135 698 137
rect 636 124 640 134
rect 646 133 650 135
rect 658 134 698 135
rect 646 131 647 133
rect 649 131 650 133
rect 646 130 650 131
rect 636 122 637 124
rect 639 122 640 124
rect 636 120 640 122
rect 643 126 650 130
rect 643 115 647 126
rect 686 121 690 126
rect 686 119 687 121
rect 689 119 690 121
rect 629 114 647 115
rect 629 112 631 114
rect 633 113 647 114
rect 633 112 658 113
rect 629 111 654 112
rect 643 110 654 111
rect 656 110 658 112
rect 643 109 658 110
rect 663 112 667 114
rect 663 110 664 112
rect 666 110 667 112
rect 663 105 667 110
rect 686 117 690 119
rect 694 123 698 134
rect 694 121 700 123
rect 694 119 697 121
rect 699 119 700 121
rect 694 117 700 119
rect 694 114 698 117
rect 678 110 698 114
rect 678 106 682 110
rect 642 104 664 105
rect 633 101 637 103
rect 642 102 644 104
rect 646 103 664 104
rect 666 103 667 105
rect 646 102 667 103
rect 672 105 682 106
rect 672 103 674 105
rect 676 103 682 105
rect 672 102 682 103
rect 733 138 737 142
rect 756 138 780 142
rect 720 137 760 138
rect 720 135 734 137
rect 736 135 760 137
rect 720 134 760 135
rect 720 123 724 134
rect 768 133 772 135
rect 776 134 782 138
rect 768 131 769 133
rect 771 131 772 133
rect 768 130 772 131
rect 768 126 775 130
rect 718 121 724 123
rect 718 119 719 121
rect 721 119 724 121
rect 718 117 724 119
rect 728 121 732 126
rect 728 119 729 121
rect 731 119 732 121
rect 728 117 732 119
rect 720 114 724 117
rect 720 110 740 114
rect 736 106 740 110
rect 771 115 775 126
rect 778 124 782 134
rect 778 122 779 124
rect 781 122 782 124
rect 778 120 782 122
rect 771 114 789 115
rect 751 112 755 114
rect 771 113 785 114
rect 751 110 752 112
rect 754 110 755 112
rect 736 105 746 106
rect 736 103 742 105
rect 744 103 746 105
rect 736 102 746 103
rect 751 105 755 110
rect 760 112 785 113
rect 787 112 789 114
rect 760 110 762 112
rect 764 111 789 112
rect 764 110 775 111
rect 760 109 775 110
rect 814 138 818 142
rect 814 134 829 138
rect 804 125 810 126
rect 825 121 829 134
rect 832 131 833 142
rect 825 119 826 121
rect 828 119 829 121
rect 825 113 829 119
rect 860 138 864 143
rect 869 143 875 152
rect 900 150 902 152
rect 904 150 906 152
rect 900 149 906 150
rect 935 150 937 152
rect 939 150 941 152
rect 869 141 871 143
rect 873 141 875 143
rect 935 145 941 150
rect 957 150 959 152
rect 961 150 963 152
rect 935 143 937 145
rect 939 143 941 145
rect 935 142 941 143
rect 948 144 952 146
rect 948 142 949 144
rect 951 142 952 144
rect 957 145 963 150
rect 957 143 959 145
rect 961 143 963 145
rect 957 142 963 143
rect 989 150 991 152
rect 993 150 995 152
rect 989 145 995 150
rect 1011 150 1013 152
rect 1015 150 1017 152
rect 989 143 991 145
rect 993 143 995 145
rect 989 142 995 143
rect 1000 144 1004 146
rect 1000 142 1001 144
rect 1003 142 1004 144
rect 1011 145 1017 150
rect 1046 150 1048 152
rect 1050 150 1052 152
rect 1046 149 1052 150
rect 1087 150 1089 152
rect 1091 150 1093 152
rect 1087 149 1093 150
rect 1011 143 1013 145
rect 1015 143 1017 145
rect 1011 142 1017 143
rect 1068 145 1085 146
rect 1068 143 1070 145
rect 1072 143 1085 145
rect 1068 142 1085 143
rect 1116 145 1122 152
rect 1116 143 1118 145
rect 1120 143 1122 145
rect 1116 142 1122 143
rect 1127 145 1131 147
rect 1127 143 1128 145
rect 1130 143 1131 145
rect 869 140 875 141
rect 860 136 861 138
rect 863 137 864 138
rect 863 136 877 137
rect 860 133 877 136
rect 811 112 829 113
rect 811 110 813 112
rect 815 110 829 112
rect 811 109 829 110
rect 873 121 877 133
rect 873 119 874 121
rect 876 119 877 121
rect 873 114 877 119
rect 865 110 877 114
rect 865 106 869 110
rect 880 107 881 109
rect 751 103 752 105
rect 754 104 776 105
rect 754 103 772 104
rect 751 102 772 103
rect 774 102 776 104
rect 642 101 667 102
rect 751 101 776 102
rect 781 101 785 103
rect 849 105 869 106
rect 849 103 851 105
rect 853 103 869 105
rect 849 102 869 103
rect 905 138 929 142
rect 948 138 952 142
rect 903 134 909 138
rect 925 137 965 138
rect 925 135 949 137
rect 951 135 965 137
rect 903 124 907 134
rect 913 133 917 135
rect 925 134 965 135
rect 913 131 914 133
rect 916 131 917 133
rect 913 130 917 131
rect 903 122 904 124
rect 906 122 907 124
rect 903 120 907 122
rect 910 126 917 130
rect 910 115 914 126
rect 953 121 957 126
rect 953 119 954 121
rect 956 119 957 121
rect 896 114 914 115
rect 896 112 898 114
rect 900 113 914 114
rect 900 112 925 113
rect 896 111 921 112
rect 910 110 921 111
rect 923 110 925 112
rect 910 109 925 110
rect 930 112 934 114
rect 930 110 931 112
rect 933 110 934 112
rect 930 105 934 110
rect 953 117 957 119
rect 961 123 965 134
rect 961 121 967 123
rect 961 119 964 121
rect 966 119 967 121
rect 961 117 967 119
rect 961 114 965 117
rect 945 110 965 114
rect 945 106 949 110
rect 909 104 931 105
rect 900 101 904 103
rect 909 102 911 104
rect 913 103 931 104
rect 933 103 934 105
rect 913 102 934 103
rect 939 105 949 106
rect 939 103 941 105
rect 943 103 949 105
rect 939 102 949 103
rect 1000 138 1004 142
rect 1023 138 1047 142
rect 987 137 1027 138
rect 987 135 1001 137
rect 1003 135 1027 137
rect 987 134 1027 135
rect 987 123 991 134
rect 1035 133 1039 135
rect 1043 134 1049 138
rect 1035 131 1036 133
rect 1038 131 1039 133
rect 1035 130 1039 131
rect 1035 126 1042 130
rect 985 121 991 123
rect 985 119 986 121
rect 988 119 991 121
rect 985 117 991 119
rect 995 121 999 126
rect 995 119 996 121
rect 998 119 999 121
rect 995 117 999 119
rect 987 114 991 117
rect 987 110 1007 114
rect 1003 106 1007 110
rect 1038 115 1042 126
rect 1045 124 1049 134
rect 1045 122 1046 124
rect 1048 122 1049 124
rect 1045 120 1049 122
rect 1038 114 1056 115
rect 1018 112 1022 114
rect 1038 113 1052 114
rect 1018 110 1019 112
rect 1021 110 1022 112
rect 1003 105 1013 106
rect 1003 103 1009 105
rect 1011 103 1013 105
rect 1003 102 1013 103
rect 1018 105 1022 110
rect 1027 112 1052 113
rect 1054 112 1056 114
rect 1027 110 1029 112
rect 1031 111 1056 112
rect 1031 110 1042 111
rect 1027 109 1042 110
rect 1081 138 1085 142
rect 1081 134 1096 138
rect 1071 125 1077 126
rect 1092 121 1096 134
rect 1099 131 1100 142
rect 1092 119 1093 121
rect 1095 119 1096 121
rect 1092 113 1096 119
rect 1127 138 1131 143
rect 1136 143 1142 152
rect 1167 150 1169 152
rect 1171 150 1173 152
rect 1167 149 1173 150
rect 1202 150 1204 152
rect 1206 150 1208 152
rect 1136 141 1138 143
rect 1140 141 1142 143
rect 1202 145 1208 150
rect 1224 150 1226 152
rect 1228 150 1230 152
rect 1202 143 1204 145
rect 1206 143 1208 145
rect 1202 142 1208 143
rect 1215 144 1219 146
rect 1215 142 1216 144
rect 1218 142 1219 144
rect 1224 145 1230 150
rect 1224 143 1226 145
rect 1228 143 1230 145
rect 1224 142 1230 143
rect 1256 150 1258 152
rect 1260 150 1262 152
rect 1256 145 1262 150
rect 1278 150 1280 152
rect 1282 150 1284 152
rect 1256 143 1258 145
rect 1260 143 1262 145
rect 1256 142 1262 143
rect 1267 144 1271 146
rect 1267 142 1268 144
rect 1270 142 1271 144
rect 1278 145 1284 150
rect 1313 150 1315 152
rect 1317 150 1319 152
rect 1313 149 1319 150
rect 1354 150 1356 152
rect 1358 150 1360 152
rect 1354 149 1360 150
rect 1278 143 1280 145
rect 1282 143 1284 145
rect 1278 142 1284 143
rect 1335 145 1352 146
rect 1335 143 1337 145
rect 1339 143 1352 145
rect 1335 142 1352 143
rect 1383 145 1389 152
rect 1383 143 1385 145
rect 1387 143 1389 145
rect 1383 142 1389 143
rect 1394 145 1398 147
rect 1394 143 1395 145
rect 1397 143 1398 145
rect 1136 140 1142 141
rect 1127 136 1128 138
rect 1130 137 1131 138
rect 1130 136 1144 137
rect 1127 133 1144 136
rect 1078 112 1096 113
rect 1078 110 1080 112
rect 1082 110 1096 112
rect 1078 109 1096 110
rect 1140 121 1144 133
rect 1140 119 1141 121
rect 1143 119 1144 121
rect 1140 114 1144 119
rect 1132 110 1144 114
rect 1132 106 1136 110
rect 1147 107 1148 109
rect 1018 103 1019 105
rect 1021 104 1043 105
rect 1021 103 1039 104
rect 1018 102 1039 103
rect 1041 102 1043 104
rect 909 101 934 102
rect 1018 101 1043 102
rect 1048 101 1052 103
rect 1116 105 1136 106
rect 1116 103 1118 105
rect 1120 103 1136 105
rect 1116 102 1136 103
rect 1172 138 1196 142
rect 1215 138 1219 142
rect 1170 134 1176 138
rect 1192 137 1232 138
rect 1192 135 1216 137
rect 1218 135 1232 137
rect 1170 124 1174 134
rect 1180 133 1184 135
rect 1192 134 1232 135
rect 1180 131 1181 133
rect 1183 131 1184 133
rect 1180 130 1184 131
rect 1170 122 1171 124
rect 1173 122 1174 124
rect 1170 120 1174 122
rect 1177 126 1184 130
rect 1177 115 1181 126
rect 1220 121 1224 126
rect 1220 119 1221 121
rect 1223 119 1224 121
rect 1163 114 1181 115
rect 1163 112 1165 114
rect 1167 113 1181 114
rect 1167 112 1192 113
rect 1163 111 1188 112
rect 1177 110 1188 111
rect 1190 110 1192 112
rect 1177 109 1192 110
rect 1197 112 1201 114
rect 1197 110 1198 112
rect 1200 110 1201 112
rect 1197 105 1201 110
rect 1220 117 1224 119
rect 1228 123 1232 134
rect 1228 121 1234 123
rect 1228 119 1231 121
rect 1233 119 1234 121
rect 1228 117 1234 119
rect 1228 114 1232 117
rect 1212 110 1232 114
rect 1212 106 1216 110
rect 1176 104 1198 105
rect 1167 101 1171 103
rect 1176 102 1178 104
rect 1180 103 1198 104
rect 1200 103 1201 105
rect 1180 102 1201 103
rect 1206 105 1216 106
rect 1206 103 1208 105
rect 1210 103 1216 105
rect 1206 102 1216 103
rect 1267 138 1271 142
rect 1290 138 1314 142
rect 1254 137 1294 138
rect 1254 135 1268 137
rect 1270 135 1294 137
rect 1254 134 1294 135
rect 1254 123 1258 134
rect 1302 133 1306 135
rect 1310 134 1316 138
rect 1302 131 1303 133
rect 1305 131 1306 133
rect 1302 130 1306 131
rect 1302 126 1309 130
rect 1252 121 1258 123
rect 1252 119 1253 121
rect 1255 119 1258 121
rect 1252 117 1258 119
rect 1262 121 1266 126
rect 1262 119 1263 121
rect 1265 119 1266 121
rect 1262 117 1266 119
rect 1254 114 1258 117
rect 1254 110 1274 114
rect 1270 106 1274 110
rect 1305 115 1309 126
rect 1312 124 1316 134
rect 1312 122 1313 124
rect 1315 122 1316 124
rect 1312 120 1316 122
rect 1305 114 1323 115
rect 1285 112 1289 114
rect 1305 113 1319 114
rect 1285 110 1286 112
rect 1288 110 1289 112
rect 1270 105 1280 106
rect 1270 103 1276 105
rect 1278 103 1280 105
rect 1270 102 1280 103
rect 1285 105 1289 110
rect 1294 112 1319 113
rect 1321 112 1323 114
rect 1294 110 1296 112
rect 1298 111 1323 112
rect 1298 110 1309 111
rect 1294 109 1309 110
rect 1348 138 1352 142
rect 1348 134 1363 138
rect 1338 125 1344 126
rect 1359 121 1363 134
rect 1366 131 1367 142
rect 1359 119 1360 121
rect 1362 119 1363 121
rect 1359 113 1363 119
rect 1394 138 1398 143
rect 1403 143 1409 152
rect 1434 150 1436 152
rect 1438 150 1440 152
rect 1434 149 1440 150
rect 1469 150 1471 152
rect 1473 150 1475 152
rect 1403 141 1405 143
rect 1407 141 1409 143
rect 1469 145 1475 150
rect 1491 150 1493 152
rect 1495 150 1497 152
rect 1469 143 1471 145
rect 1473 143 1475 145
rect 1469 142 1475 143
rect 1482 144 1486 146
rect 1482 142 1483 144
rect 1485 142 1486 144
rect 1491 145 1497 150
rect 1491 143 1493 145
rect 1495 143 1497 145
rect 1491 142 1497 143
rect 1523 150 1525 152
rect 1527 150 1529 152
rect 1523 145 1529 150
rect 1545 150 1547 152
rect 1549 150 1551 152
rect 1523 143 1525 145
rect 1527 143 1529 145
rect 1523 142 1529 143
rect 1534 144 1538 146
rect 1534 142 1535 144
rect 1537 142 1538 144
rect 1545 145 1551 150
rect 1580 150 1582 152
rect 1584 150 1586 152
rect 1580 149 1586 150
rect 1621 150 1623 152
rect 1625 150 1627 152
rect 1621 149 1627 150
rect 1545 143 1547 145
rect 1549 143 1551 145
rect 1545 142 1551 143
rect 1602 145 1619 146
rect 1602 143 1604 145
rect 1606 143 1619 145
rect 1602 142 1619 143
rect 1650 145 1656 152
rect 1650 143 1652 145
rect 1654 143 1656 145
rect 1650 142 1656 143
rect 1661 145 1665 147
rect 1661 143 1662 145
rect 1664 143 1665 145
rect 1403 140 1409 141
rect 1394 136 1395 138
rect 1397 137 1398 138
rect 1397 136 1411 137
rect 1394 133 1411 136
rect 1345 112 1363 113
rect 1345 110 1347 112
rect 1349 110 1363 112
rect 1345 109 1363 110
rect 1407 121 1411 133
rect 1407 119 1408 121
rect 1410 119 1411 121
rect 1407 114 1411 119
rect 1399 110 1411 114
rect 1399 106 1403 110
rect 1414 107 1415 109
rect 1285 103 1286 105
rect 1288 104 1310 105
rect 1288 103 1306 104
rect 1285 102 1306 103
rect 1308 102 1310 104
rect 1176 101 1201 102
rect 1285 101 1310 102
rect 1315 101 1319 103
rect 1383 105 1403 106
rect 1383 103 1385 105
rect 1387 103 1403 105
rect 1383 102 1403 103
rect 1439 138 1463 142
rect 1482 138 1486 142
rect 1437 134 1443 138
rect 1459 137 1499 138
rect 1459 135 1483 137
rect 1485 135 1499 137
rect 1437 124 1441 134
rect 1447 133 1451 135
rect 1459 134 1499 135
rect 1447 131 1448 133
rect 1450 131 1451 133
rect 1447 130 1451 131
rect 1437 122 1438 124
rect 1440 122 1441 124
rect 1437 120 1441 122
rect 1444 126 1451 130
rect 1444 115 1448 126
rect 1487 121 1491 126
rect 1487 119 1488 121
rect 1490 119 1491 121
rect 1430 114 1448 115
rect 1430 112 1432 114
rect 1434 113 1448 114
rect 1434 112 1459 113
rect 1430 111 1455 112
rect 1444 110 1455 111
rect 1457 110 1459 112
rect 1444 109 1459 110
rect 1464 112 1468 114
rect 1464 110 1465 112
rect 1467 110 1468 112
rect 1464 105 1468 110
rect 1487 117 1491 119
rect 1495 123 1499 134
rect 1495 121 1501 123
rect 1495 119 1498 121
rect 1500 119 1501 121
rect 1495 117 1501 119
rect 1495 114 1499 117
rect 1479 110 1499 114
rect 1479 106 1483 110
rect 1443 104 1465 105
rect 1434 101 1438 103
rect 1443 102 1445 104
rect 1447 103 1465 104
rect 1467 103 1468 105
rect 1447 102 1468 103
rect 1473 105 1483 106
rect 1473 103 1475 105
rect 1477 103 1483 105
rect 1473 102 1483 103
rect 1534 138 1538 142
rect 1557 138 1581 142
rect 1521 137 1561 138
rect 1521 135 1535 137
rect 1537 135 1561 137
rect 1521 134 1561 135
rect 1521 123 1525 134
rect 1569 133 1573 135
rect 1577 134 1583 138
rect 1569 131 1570 133
rect 1572 131 1573 133
rect 1569 130 1573 131
rect 1569 126 1576 130
rect 1519 121 1525 123
rect 1519 119 1520 121
rect 1522 119 1525 121
rect 1519 117 1525 119
rect 1529 121 1533 126
rect 1529 119 1530 121
rect 1532 119 1533 121
rect 1529 117 1533 119
rect 1521 114 1525 117
rect 1521 110 1541 114
rect 1537 106 1541 110
rect 1572 115 1576 126
rect 1579 124 1583 134
rect 1579 122 1580 124
rect 1582 122 1583 124
rect 1579 120 1583 122
rect 1572 114 1590 115
rect 1552 112 1556 114
rect 1572 113 1586 114
rect 1552 110 1553 112
rect 1555 110 1556 112
rect 1537 105 1547 106
rect 1537 103 1543 105
rect 1545 103 1547 105
rect 1537 102 1547 103
rect 1552 105 1556 110
rect 1561 112 1586 113
rect 1588 112 1590 114
rect 1561 110 1563 112
rect 1565 111 1590 112
rect 1565 110 1576 111
rect 1561 109 1576 110
rect 1615 138 1619 142
rect 1615 134 1630 138
rect 1605 125 1611 126
rect 1626 121 1630 134
rect 1633 131 1634 142
rect 1626 119 1627 121
rect 1629 119 1630 121
rect 1626 113 1630 119
rect 1661 138 1665 143
rect 1670 143 1676 152
rect 1701 150 1703 152
rect 1705 150 1707 152
rect 1701 149 1707 150
rect 1736 150 1738 152
rect 1740 150 1742 152
rect 1670 141 1672 143
rect 1674 141 1676 143
rect 1736 145 1742 150
rect 1758 150 1760 152
rect 1762 150 1764 152
rect 1736 143 1738 145
rect 1740 143 1742 145
rect 1736 142 1742 143
rect 1749 144 1753 146
rect 1749 142 1750 144
rect 1752 142 1753 144
rect 1758 145 1764 150
rect 1758 143 1760 145
rect 1762 143 1764 145
rect 1758 142 1764 143
rect 1790 150 1792 152
rect 1794 150 1796 152
rect 1790 145 1796 150
rect 1812 150 1814 152
rect 1816 150 1818 152
rect 1790 143 1792 145
rect 1794 143 1796 145
rect 1790 142 1796 143
rect 1801 144 1805 146
rect 1801 142 1802 144
rect 1804 142 1805 144
rect 1812 145 1818 150
rect 1847 150 1849 152
rect 1851 150 1853 152
rect 1847 149 1853 150
rect 1888 150 1890 152
rect 1892 150 1894 152
rect 1888 149 1894 150
rect 1931 150 1932 152
rect 1934 150 1935 152
rect 1812 143 1814 145
rect 1816 143 1818 145
rect 1812 142 1818 143
rect 1869 145 1886 146
rect 1869 143 1871 145
rect 1873 143 1886 145
rect 1869 142 1886 143
rect 1670 140 1676 141
rect 1661 136 1662 138
rect 1664 137 1665 138
rect 1664 136 1678 137
rect 1661 133 1678 136
rect 1612 112 1630 113
rect 1612 110 1614 112
rect 1616 110 1630 112
rect 1612 109 1630 110
rect 1674 121 1678 133
rect 1674 119 1675 121
rect 1677 119 1678 121
rect 1674 114 1678 119
rect 1666 110 1678 114
rect 1666 106 1670 110
rect 1681 107 1682 109
rect 1552 103 1553 105
rect 1555 104 1577 105
rect 1555 103 1573 104
rect 1552 102 1573 103
rect 1575 102 1577 104
rect 1443 101 1468 102
rect 1552 101 1577 102
rect 1582 101 1586 103
rect 1650 105 1670 106
rect 1650 103 1652 105
rect 1654 103 1670 105
rect 1650 102 1670 103
rect 1706 138 1730 142
rect 1749 138 1753 142
rect 1704 134 1710 138
rect 1726 137 1766 138
rect 1726 135 1750 137
rect 1752 135 1766 137
rect 1704 124 1708 134
rect 1714 133 1718 135
rect 1726 134 1766 135
rect 1714 131 1715 133
rect 1717 131 1718 133
rect 1714 130 1718 131
rect 1704 122 1705 124
rect 1707 122 1708 124
rect 1704 120 1708 122
rect 1711 126 1718 130
rect 1711 115 1715 126
rect 1754 121 1758 126
rect 1754 119 1755 121
rect 1757 119 1758 121
rect 1697 114 1715 115
rect 1697 112 1699 114
rect 1701 113 1715 114
rect 1701 112 1726 113
rect 1697 111 1722 112
rect 1711 110 1722 111
rect 1724 110 1726 112
rect 1711 109 1726 110
rect 1731 112 1735 114
rect 1731 110 1732 112
rect 1734 110 1735 112
rect 1731 105 1735 110
rect 1754 117 1758 119
rect 1762 123 1766 134
rect 1762 121 1768 123
rect 1762 119 1765 121
rect 1767 119 1768 121
rect 1762 117 1768 119
rect 1762 114 1766 117
rect 1746 110 1766 114
rect 1746 106 1750 110
rect 1710 104 1732 105
rect 1701 101 1705 103
rect 1710 102 1712 104
rect 1714 103 1732 104
rect 1734 103 1735 105
rect 1714 102 1735 103
rect 1740 105 1750 106
rect 1740 103 1742 105
rect 1744 103 1750 105
rect 1740 102 1750 103
rect 1801 138 1805 142
rect 1824 138 1848 142
rect 1788 137 1828 138
rect 1788 135 1802 137
rect 1804 135 1828 137
rect 1788 134 1828 135
rect 1788 123 1792 134
rect 1836 133 1840 135
rect 1844 134 1850 138
rect 1836 131 1837 133
rect 1839 131 1840 133
rect 1836 130 1840 131
rect 1836 126 1843 130
rect 1786 121 1792 123
rect 1786 119 1787 121
rect 1789 119 1792 121
rect 1786 117 1792 119
rect 1796 121 1800 126
rect 1796 119 1797 121
rect 1799 119 1800 121
rect 1796 117 1800 119
rect 1788 114 1792 117
rect 1788 110 1808 114
rect 1804 106 1808 110
rect 1839 115 1843 126
rect 1846 124 1850 134
rect 1846 122 1847 124
rect 1849 122 1850 124
rect 1846 120 1850 122
rect 1839 114 1857 115
rect 1819 112 1823 114
rect 1839 113 1853 114
rect 1819 110 1820 112
rect 1822 110 1823 112
rect 1804 105 1814 106
rect 1804 103 1810 105
rect 1812 103 1814 105
rect 1804 102 1814 103
rect 1819 105 1823 110
rect 1828 112 1853 113
rect 1855 112 1857 114
rect 1828 110 1830 112
rect 1832 111 1857 112
rect 1882 138 1886 142
rect 1882 134 1897 138
rect 1872 125 1878 126
rect 1893 121 1897 134
rect 1900 131 1901 142
rect 1893 119 1894 121
rect 1896 119 1897 121
rect 1893 113 1897 119
rect 1931 145 1935 150
rect 1987 150 1989 152
rect 1991 150 1993 152
rect 1987 149 1993 150
rect 2022 150 2024 152
rect 2026 150 2028 152
rect 1931 143 1932 145
rect 1934 143 1935 145
rect 1931 141 1935 143
rect 1939 146 1972 147
rect 1939 144 1968 146
rect 1970 144 1972 146
rect 1939 143 1972 144
rect 2022 145 2028 150
rect 2044 150 2046 152
rect 2048 150 2050 152
rect 2022 143 2024 145
rect 2026 143 2028 145
rect 1939 132 1943 143
rect 2022 142 2028 143
rect 2035 144 2039 146
rect 2035 142 2036 144
rect 2038 142 2039 144
rect 2044 145 2050 150
rect 2044 143 2046 145
rect 2048 143 2050 145
rect 2044 142 2050 143
rect 2076 150 2078 152
rect 2080 150 2082 152
rect 2076 145 2082 150
rect 2098 150 2100 152
rect 2102 150 2104 152
rect 2076 143 2078 145
rect 2080 143 2082 145
rect 2076 142 2082 143
rect 2087 144 2091 146
rect 2087 142 2088 144
rect 2090 142 2091 144
rect 2098 145 2104 150
rect 2133 150 2135 152
rect 2137 150 2139 152
rect 2133 149 2139 150
rect 2174 150 2176 152
rect 2178 150 2180 152
rect 2174 149 2180 150
rect 2210 150 2211 152
rect 2213 150 2214 152
rect 2210 148 2214 150
rect 2243 150 2245 152
rect 2247 150 2249 152
rect 2243 149 2249 150
rect 2278 150 2279 152
rect 2281 150 2282 152
rect 2278 148 2282 150
rect 2311 150 2313 152
rect 2315 150 2317 152
rect 2311 149 2317 150
rect 2098 143 2100 145
rect 2102 143 2104 145
rect 2098 142 2104 143
rect 2155 145 2172 146
rect 2155 143 2157 145
rect 2159 143 2172 145
rect 2155 142 2172 143
rect 1920 131 1943 132
rect 1920 129 1922 131
rect 1924 129 1943 131
rect 1920 128 1943 129
rect 1920 122 1924 128
rect 1832 110 1843 111
rect 1828 109 1843 110
rect 1879 112 1897 113
rect 1879 110 1881 112
rect 1883 110 1897 112
rect 1879 109 1897 110
rect 1913 118 1924 122
rect 1913 112 1917 118
rect 1939 122 1943 128
rect 1947 138 1951 140
rect 1947 136 1948 138
rect 1950 136 1951 138
rect 1947 131 1951 136
rect 1947 129 1948 131
rect 1950 130 1951 131
rect 1950 129 1963 130
rect 1947 126 1963 129
rect 1959 124 1963 126
rect 1959 122 1964 124
rect 1939 121 1955 122
rect 1939 119 1951 121
rect 1953 119 1955 121
rect 1939 118 1955 119
rect 1959 120 1961 122
rect 1963 120 1964 122
rect 1959 118 1964 120
rect 1913 110 1914 112
rect 1916 110 1917 112
rect 1913 108 1917 110
rect 1959 114 1963 118
rect 1939 110 1963 114
rect 1939 107 1943 110
rect 1939 105 1940 107
rect 1942 105 1943 107
rect 1819 103 1820 105
rect 1822 104 1844 105
rect 1822 103 1840 104
rect 1819 102 1840 103
rect 1842 102 1844 104
rect 1710 101 1735 102
rect 1819 101 1844 102
rect 1849 101 1853 103
rect 1926 104 1932 105
rect 1926 102 1928 104
rect 1930 102 1932 104
rect 1939 103 1943 105
rect 1992 138 2016 142
rect 2035 138 2039 142
rect 1990 134 1996 138
rect 2012 137 2052 138
rect 2012 135 2036 137
rect 2038 135 2052 137
rect 1990 124 1994 134
rect 2000 133 2004 135
rect 2012 134 2052 135
rect 2000 131 2001 133
rect 2003 131 2004 133
rect 2000 130 2004 131
rect 1990 122 1991 124
rect 1993 122 1994 124
rect 1990 120 1994 122
rect 1997 126 2004 130
rect 1997 115 2001 126
rect 2040 121 2044 126
rect 2040 119 2041 121
rect 2043 119 2044 121
rect 1983 114 2001 115
rect 1983 112 1985 114
rect 1987 113 2001 114
rect 1987 112 2012 113
rect 1983 111 2008 112
rect 1997 110 2008 111
rect 2010 110 2012 112
rect 1997 109 2012 110
rect 2017 112 2021 114
rect 2017 110 2018 112
rect 2020 110 2021 112
rect 2017 105 2021 110
rect 2040 117 2044 119
rect 2048 123 2052 134
rect 2048 121 2054 123
rect 2048 119 2051 121
rect 2053 119 2054 121
rect 2048 117 2054 119
rect 2048 114 2052 117
rect 2032 110 2052 114
rect 2032 106 2036 110
rect 1996 104 2018 105
rect 99 99 100 101
rect 102 99 103 101
rect 247 99 248 101
rect 250 99 251 101
rect 99 96 103 99
rect 155 98 161 99
rect 155 96 157 98
rect 159 96 161 98
rect 189 98 195 99
rect 189 96 191 98
rect 193 96 195 98
rect 247 96 251 99
rect 267 99 273 100
rect 267 97 269 99
rect 271 97 273 99
rect 267 96 273 97
rect 286 99 292 100
rect 286 97 288 99
rect 290 97 292 99
rect 286 96 292 97
rect 366 99 367 101
rect 369 99 370 101
rect 514 99 515 101
rect 517 99 518 101
rect 366 96 370 99
rect 422 98 428 99
rect 422 96 424 98
rect 426 96 428 98
rect 456 98 462 99
rect 456 96 458 98
rect 460 96 462 98
rect 514 96 518 99
rect 534 99 540 100
rect 534 97 536 99
rect 538 97 540 99
rect 534 96 540 97
rect 553 99 559 100
rect 553 97 555 99
rect 557 97 559 99
rect 553 96 559 97
rect 633 99 634 101
rect 636 99 637 101
rect 781 99 782 101
rect 784 99 785 101
rect 633 96 637 99
rect 689 98 695 99
rect 689 96 691 98
rect 693 96 695 98
rect 723 98 729 99
rect 723 96 725 98
rect 727 96 729 98
rect 781 96 785 99
rect 801 99 807 100
rect 801 97 803 99
rect 805 97 807 99
rect 801 96 807 97
rect 820 99 826 100
rect 820 97 822 99
rect 824 97 826 99
rect 820 96 826 97
rect 900 99 901 101
rect 903 99 904 101
rect 1048 99 1049 101
rect 1051 99 1052 101
rect 900 96 904 99
rect 956 98 962 99
rect 956 96 958 98
rect 960 96 962 98
rect 990 98 996 99
rect 990 96 992 98
rect 994 96 996 98
rect 1048 96 1052 99
rect 1068 99 1074 100
rect 1068 97 1070 99
rect 1072 97 1074 99
rect 1068 96 1074 97
rect 1087 99 1093 100
rect 1087 97 1089 99
rect 1091 97 1093 99
rect 1087 96 1093 97
rect 1167 99 1168 101
rect 1170 99 1171 101
rect 1315 99 1316 101
rect 1318 99 1319 101
rect 1167 96 1171 99
rect 1223 98 1229 99
rect 1223 96 1225 98
rect 1227 96 1229 98
rect 1257 98 1263 99
rect 1257 96 1259 98
rect 1261 96 1263 98
rect 1315 96 1319 99
rect 1335 99 1341 100
rect 1335 97 1337 99
rect 1339 97 1341 99
rect 1335 96 1341 97
rect 1354 99 1360 100
rect 1354 97 1356 99
rect 1358 97 1360 99
rect 1354 96 1360 97
rect 1434 99 1435 101
rect 1437 99 1438 101
rect 1582 99 1583 101
rect 1585 99 1586 101
rect 1434 96 1438 99
rect 1490 98 1496 99
rect 1490 96 1492 98
rect 1494 96 1496 98
rect 1524 98 1530 99
rect 1524 96 1526 98
rect 1528 96 1530 98
rect 1582 96 1586 99
rect 1602 99 1608 100
rect 1602 97 1604 99
rect 1606 97 1608 99
rect 1602 96 1608 97
rect 1621 99 1627 100
rect 1621 97 1623 99
rect 1625 97 1627 99
rect 1621 96 1627 97
rect 1701 99 1702 101
rect 1704 99 1705 101
rect 1849 99 1850 101
rect 1852 99 1853 101
rect 1701 96 1705 99
rect 1757 98 1763 99
rect 1757 96 1759 98
rect 1761 96 1763 98
rect 1791 98 1797 99
rect 1791 96 1793 98
rect 1795 96 1797 98
rect 1849 96 1853 99
rect 1869 99 1875 100
rect 1869 97 1871 99
rect 1873 97 1875 99
rect 1869 96 1875 97
rect 1888 99 1894 100
rect 1888 97 1890 99
rect 1892 97 1894 99
rect 1888 96 1894 97
rect 1926 96 1932 102
rect 1987 101 1991 103
rect 1996 102 1998 104
rect 2000 103 2018 104
rect 2020 103 2021 105
rect 2000 102 2021 103
rect 2026 105 2036 106
rect 2026 103 2028 105
rect 2030 103 2036 105
rect 2026 102 2036 103
rect 2087 138 2091 142
rect 2110 138 2134 142
rect 2074 137 2114 138
rect 2074 135 2088 137
rect 2090 135 2114 137
rect 2074 134 2114 135
rect 2074 123 2078 134
rect 2122 133 2126 135
rect 2130 134 2136 138
rect 2122 131 2123 133
rect 2125 131 2126 133
rect 2122 130 2126 131
rect 2122 126 2129 130
rect 2072 121 2078 123
rect 2072 119 2073 121
rect 2075 119 2078 121
rect 2072 117 2078 119
rect 2082 121 2086 126
rect 2082 119 2083 121
rect 2085 119 2086 121
rect 2082 117 2086 119
rect 2074 114 2078 117
rect 2074 110 2094 114
rect 2090 106 2094 110
rect 2125 115 2129 126
rect 2132 124 2136 134
rect 2132 122 2133 124
rect 2135 122 2136 124
rect 2132 120 2136 122
rect 2125 114 2143 115
rect 2105 112 2109 114
rect 2125 113 2139 114
rect 2105 110 2106 112
rect 2108 110 2109 112
rect 2090 105 2100 106
rect 2090 103 2096 105
rect 2098 103 2100 105
rect 2090 102 2100 103
rect 2105 105 2109 110
rect 2114 112 2139 113
rect 2141 112 2143 114
rect 2114 110 2116 112
rect 2118 111 2143 112
rect 2168 138 2172 142
rect 2168 134 2183 138
rect 2158 125 2164 126
rect 2118 110 2129 111
rect 2114 109 2129 110
rect 2179 121 2183 134
rect 2186 131 2187 142
rect 2226 142 2239 143
rect 2226 140 2228 142
rect 2230 140 2239 142
rect 2226 139 2239 140
rect 2235 135 2251 139
rect 2179 119 2180 121
rect 2182 119 2183 121
rect 2179 113 2183 119
rect 2223 131 2227 133
rect 2165 112 2183 113
rect 2165 110 2167 112
rect 2169 110 2183 112
rect 2165 109 2183 110
rect 2199 130 2224 131
rect 2199 128 2201 130
rect 2203 129 2224 130
rect 2226 129 2227 131
rect 2203 128 2227 129
rect 2199 127 2227 128
rect 2105 103 2106 105
rect 2108 104 2130 105
rect 2108 103 2126 104
rect 2105 102 2126 103
rect 2128 102 2130 104
rect 2199 107 2203 127
rect 2223 117 2227 127
rect 2243 122 2244 128
rect 2247 118 2251 135
rect 2223 115 2234 117
rect 2223 113 2231 115
rect 2233 113 2234 115
rect 2247 116 2252 118
rect 2247 114 2249 116
rect 2251 114 2252 116
rect 2223 111 2234 113
rect 2237 112 2252 114
rect 2237 110 2251 112
rect 2199 106 2205 107
rect 2199 104 2201 106
rect 2203 104 2205 106
rect 2199 103 2205 104
rect 2209 106 2215 107
rect 2209 104 2211 106
rect 2213 104 2215 106
rect 2237 105 2241 110
rect 2294 142 2307 143
rect 2294 140 2296 142
rect 2298 140 2307 142
rect 2294 139 2307 140
rect 2303 135 2319 139
rect 2291 131 2295 133
rect 1996 101 2021 102
rect 2105 101 2130 102
rect 2135 101 2139 103
rect 1987 99 1988 101
rect 1990 99 1991 101
rect 2135 99 2136 101
rect 2138 99 2139 101
rect 1987 96 1991 99
rect 2043 98 2049 99
rect 2043 96 2045 98
rect 2047 96 2049 98
rect 2077 98 2083 99
rect 2077 96 2079 98
rect 2081 96 2083 98
rect 2135 96 2139 99
rect 2155 99 2161 100
rect 2155 97 2157 99
rect 2159 97 2161 99
rect 2155 96 2161 97
rect 2174 99 2180 100
rect 2174 97 2176 99
rect 2178 97 2180 99
rect 2174 96 2180 97
rect 2209 96 2215 104
rect 2226 104 2241 105
rect 2226 102 2228 104
rect 2230 102 2241 104
rect 2226 101 2241 102
rect 2244 104 2248 106
rect 2244 102 2245 104
rect 2247 102 2248 104
rect 2267 130 2292 131
rect 2267 128 2269 130
rect 2271 129 2292 130
rect 2294 129 2295 131
rect 2271 128 2295 129
rect 2267 127 2295 128
rect 2267 107 2271 127
rect 2291 117 2295 127
rect 2311 122 2312 128
rect 2315 118 2319 135
rect 2291 115 2302 117
rect 2291 113 2299 115
rect 2301 113 2302 115
rect 2315 116 2320 118
rect 2315 114 2317 116
rect 2319 114 2320 116
rect 2291 111 2302 113
rect 2305 112 2320 114
rect 2305 110 2319 112
rect 2267 106 2273 107
rect 2267 104 2269 106
rect 2271 104 2273 106
rect 2267 103 2273 104
rect 2277 106 2283 107
rect 2277 104 2279 106
rect 2281 104 2283 106
rect 2305 105 2309 110
rect 2244 96 2248 102
rect 2277 96 2283 104
rect 2294 104 2309 105
rect 2294 102 2296 104
rect 2298 102 2309 104
rect 2294 101 2309 102
rect 2312 104 2316 106
rect 2312 102 2313 104
rect 2315 102 2316 104
rect 2312 96 2316 102
rect 99 77 103 80
rect 155 78 157 80
rect 159 78 161 80
rect 155 77 161 78
rect 189 78 191 80
rect 193 78 195 80
rect 189 77 195 78
rect 247 77 251 80
rect 99 75 100 77
rect 102 75 103 77
rect 247 75 248 77
rect 250 75 251 77
rect 267 79 273 80
rect 267 77 269 79
rect 271 77 273 79
rect 267 76 273 77
rect 286 79 292 80
rect 286 77 288 79
rect 290 77 292 79
rect 286 76 292 77
rect 366 77 370 80
rect 422 78 424 80
rect 426 78 428 80
rect 422 77 428 78
rect 456 78 458 80
rect 460 78 462 80
rect 456 77 462 78
rect 514 77 518 80
rect 366 75 367 77
rect 369 75 370 77
rect 514 75 515 77
rect 517 75 518 77
rect 534 79 540 80
rect 534 77 536 79
rect 538 77 540 79
rect 534 76 540 77
rect 553 79 559 80
rect 553 77 555 79
rect 557 77 559 79
rect 553 76 559 77
rect 633 77 637 80
rect 689 78 691 80
rect 693 78 695 80
rect 689 77 695 78
rect 723 78 725 80
rect 727 78 729 80
rect 723 77 729 78
rect 781 77 785 80
rect 633 75 634 77
rect 636 75 637 77
rect 781 75 782 77
rect 784 75 785 77
rect 801 79 807 80
rect 801 77 803 79
rect 805 77 807 79
rect 801 76 807 77
rect 820 79 826 80
rect 820 77 822 79
rect 824 77 826 79
rect 820 76 826 77
rect 900 77 904 80
rect 956 78 958 80
rect 960 78 962 80
rect 956 77 962 78
rect 990 78 992 80
rect 994 78 996 80
rect 990 77 996 78
rect 1048 77 1052 80
rect 900 75 901 77
rect 903 75 904 77
rect 1048 75 1049 77
rect 1051 75 1052 77
rect 1068 79 1074 80
rect 1068 77 1070 79
rect 1072 77 1074 79
rect 1068 76 1074 77
rect 1087 79 1093 80
rect 1087 77 1089 79
rect 1091 77 1093 79
rect 1087 76 1093 77
rect 1167 77 1171 80
rect 1223 78 1225 80
rect 1227 78 1229 80
rect 1223 77 1229 78
rect 1257 78 1259 80
rect 1261 78 1263 80
rect 1257 77 1263 78
rect 1315 77 1319 80
rect 1167 75 1168 77
rect 1170 75 1171 77
rect 1315 75 1316 77
rect 1318 75 1319 77
rect 1335 79 1341 80
rect 1335 77 1337 79
rect 1339 77 1341 79
rect 1335 76 1341 77
rect 1354 79 1360 80
rect 1354 77 1356 79
rect 1358 77 1360 79
rect 1354 76 1360 77
rect 1434 77 1438 80
rect 1490 78 1492 80
rect 1494 78 1496 80
rect 1490 77 1496 78
rect 1524 78 1526 80
rect 1528 78 1530 80
rect 1524 77 1530 78
rect 1582 77 1586 80
rect 1434 75 1435 77
rect 1437 75 1438 77
rect 1582 75 1583 77
rect 1585 75 1586 77
rect 1602 79 1608 80
rect 1602 77 1604 79
rect 1606 77 1608 79
rect 1602 76 1608 77
rect 1621 79 1627 80
rect 1621 77 1623 79
rect 1625 77 1627 79
rect 1621 76 1627 77
rect 1701 77 1705 80
rect 1757 78 1759 80
rect 1761 78 1763 80
rect 1757 77 1763 78
rect 1791 78 1793 80
rect 1795 78 1797 80
rect 1791 77 1797 78
rect 1849 77 1853 80
rect 1701 75 1702 77
rect 1704 75 1705 77
rect 1849 75 1850 77
rect 1852 75 1853 77
rect 1869 79 1875 80
rect 1869 77 1871 79
rect 1873 77 1875 79
rect 1869 76 1875 77
rect 1888 79 1894 80
rect 1888 77 1890 79
rect 1892 77 1894 79
rect 1888 76 1894 77
rect 8 73 28 74
rect 8 71 10 73
rect 12 71 28 73
rect 8 70 28 71
rect 24 66 28 70
rect 48 73 68 74
rect 48 71 50 73
rect 52 71 68 73
rect 48 70 68 71
rect 39 67 40 69
rect 24 62 36 66
rect 32 57 36 62
rect 32 55 33 57
rect 35 55 36 57
rect 32 43 36 55
rect 64 66 68 70
rect 79 67 80 69
rect 64 62 76 66
rect 72 57 76 62
rect 72 55 73 57
rect 75 55 76 57
rect 19 40 36 43
rect 19 38 20 40
rect 22 39 36 40
rect 22 38 23 39
rect 8 33 14 34
rect 8 31 10 33
rect 12 31 14 33
rect 8 24 14 31
rect 19 33 23 38
rect 72 43 76 55
rect 59 40 76 43
rect 59 38 60 40
rect 62 39 76 40
rect 62 38 63 39
rect 19 31 20 33
rect 22 31 23 33
rect 19 29 23 31
rect 28 35 34 36
rect 28 33 30 35
rect 32 33 34 35
rect 48 33 54 34
rect 28 24 34 33
rect 48 31 50 33
rect 52 31 54 33
rect 48 24 54 31
rect 59 33 63 38
rect 99 73 103 75
rect 108 74 133 75
rect 217 74 242 75
rect 108 72 110 74
rect 112 73 133 74
rect 112 72 130 73
rect 108 71 130 72
rect 132 71 133 73
rect 109 66 124 67
rect 109 65 120 66
rect 95 64 120 65
rect 122 64 124 66
rect 95 62 97 64
rect 99 63 124 64
rect 129 66 133 71
rect 138 73 148 74
rect 138 71 140 73
rect 142 71 148 73
rect 138 70 148 71
rect 129 64 130 66
rect 132 64 133 66
rect 99 62 113 63
rect 129 62 133 64
rect 95 61 113 62
rect 102 54 106 56
rect 102 52 103 54
rect 105 52 106 54
rect 102 42 106 52
rect 109 50 113 61
rect 144 66 148 70
rect 144 62 164 66
rect 160 59 164 62
rect 152 57 156 59
rect 152 55 153 57
rect 155 55 156 57
rect 152 50 156 55
rect 160 57 166 59
rect 160 55 163 57
rect 165 55 166 57
rect 160 53 166 55
rect 109 46 116 50
rect 112 45 116 46
rect 112 43 113 45
rect 115 43 116 45
rect 102 38 108 42
rect 112 41 116 43
rect 160 42 164 53
rect 124 41 164 42
rect 124 39 148 41
rect 150 39 164 41
rect 124 38 164 39
rect 59 31 60 33
rect 62 31 63 33
rect 59 29 63 31
rect 68 35 74 36
rect 68 33 70 35
rect 72 33 74 35
rect 104 34 128 38
rect 147 34 151 38
rect 202 73 212 74
rect 202 71 208 73
rect 210 71 212 73
rect 202 70 212 71
rect 217 73 238 74
rect 217 71 218 73
rect 220 72 238 73
rect 240 72 242 74
rect 247 73 251 75
rect 220 71 242 72
rect 202 66 206 70
rect 186 62 206 66
rect 186 59 190 62
rect 184 57 190 59
rect 184 55 185 57
rect 187 55 190 57
rect 184 53 190 55
rect 186 42 190 53
rect 194 57 198 59
rect 217 66 221 71
rect 315 73 335 74
rect 315 71 317 73
rect 319 71 335 73
rect 315 70 335 71
rect 217 64 218 66
rect 220 64 221 66
rect 217 62 221 64
rect 226 66 241 67
rect 226 64 228 66
rect 230 65 241 66
rect 230 64 255 65
rect 226 63 251 64
rect 237 62 251 63
rect 253 62 255 64
rect 237 61 255 62
rect 194 55 195 57
rect 197 55 198 57
rect 194 50 198 55
rect 237 50 241 61
rect 234 46 241 50
rect 244 54 248 56
rect 244 52 245 54
rect 247 52 248 54
rect 234 45 238 46
rect 234 43 235 45
rect 237 43 238 45
rect 186 41 226 42
rect 234 41 238 43
rect 244 42 248 52
rect 277 66 295 67
rect 277 64 279 66
rect 281 64 295 66
rect 277 63 295 64
rect 291 57 295 63
rect 291 55 292 57
rect 294 55 295 57
rect 270 50 276 51
rect 186 39 200 41
rect 202 39 226 41
rect 186 38 226 39
rect 242 38 248 42
rect 199 34 203 38
rect 222 34 246 38
rect 291 42 295 55
rect 280 38 295 42
rect 280 34 284 38
rect 298 34 299 45
rect 331 66 335 70
rect 346 67 347 69
rect 331 62 343 66
rect 339 57 343 62
rect 339 55 340 57
rect 342 55 343 57
rect 339 43 343 55
rect 326 40 343 43
rect 326 38 327 40
rect 329 39 343 40
rect 329 38 330 39
rect 68 24 74 33
rect 134 33 140 34
rect 134 31 136 33
rect 138 31 140 33
rect 99 26 105 27
rect 99 24 101 26
rect 103 24 105 26
rect 134 26 140 31
rect 147 32 148 34
rect 150 32 151 34
rect 147 30 151 32
rect 156 33 162 34
rect 156 31 158 33
rect 160 31 162 33
rect 134 24 136 26
rect 138 24 140 26
rect 156 26 162 31
rect 156 24 158 26
rect 160 24 162 26
rect 188 33 194 34
rect 188 31 190 33
rect 192 31 194 33
rect 188 26 194 31
rect 199 32 200 34
rect 202 32 203 34
rect 199 30 203 32
rect 210 33 216 34
rect 210 31 212 33
rect 214 31 216 33
rect 188 24 190 26
rect 192 24 194 26
rect 210 26 216 31
rect 267 33 284 34
rect 267 31 269 33
rect 271 31 284 33
rect 267 30 284 31
rect 315 33 321 34
rect 315 31 317 33
rect 319 31 321 33
rect 210 24 212 26
rect 214 24 216 26
rect 245 26 251 27
rect 245 24 247 26
rect 249 24 251 26
rect 286 26 292 27
rect 286 24 288 26
rect 290 24 292 26
rect 315 24 321 31
rect 326 33 330 38
rect 366 73 370 75
rect 375 74 400 75
rect 484 74 509 75
rect 375 72 377 74
rect 379 73 400 74
rect 379 72 397 73
rect 375 71 397 72
rect 399 71 400 73
rect 376 66 391 67
rect 376 65 387 66
rect 362 64 387 65
rect 389 64 391 66
rect 362 62 364 64
rect 366 63 391 64
rect 396 66 400 71
rect 405 73 415 74
rect 405 71 407 73
rect 409 71 415 73
rect 405 70 415 71
rect 396 64 397 66
rect 399 64 400 66
rect 366 62 380 63
rect 396 62 400 64
rect 362 61 380 62
rect 369 54 373 56
rect 369 52 370 54
rect 372 52 373 54
rect 369 42 373 52
rect 376 50 380 61
rect 411 66 415 70
rect 411 62 431 66
rect 427 59 431 62
rect 419 57 423 59
rect 419 55 420 57
rect 422 55 423 57
rect 419 50 423 55
rect 427 57 433 59
rect 427 55 430 57
rect 432 55 433 57
rect 427 53 433 55
rect 376 46 383 50
rect 379 45 383 46
rect 379 43 380 45
rect 382 43 383 45
rect 369 38 375 42
rect 379 41 383 43
rect 427 42 431 53
rect 391 41 431 42
rect 391 39 415 41
rect 417 39 431 41
rect 391 38 431 39
rect 326 31 327 33
rect 329 31 330 33
rect 326 29 330 31
rect 335 35 341 36
rect 335 33 337 35
rect 339 33 341 35
rect 371 34 395 38
rect 414 34 418 38
rect 469 73 479 74
rect 469 71 475 73
rect 477 71 479 73
rect 469 70 479 71
rect 484 73 505 74
rect 484 71 485 73
rect 487 72 505 73
rect 507 72 509 74
rect 514 73 518 75
rect 487 71 509 72
rect 469 66 473 70
rect 453 62 473 66
rect 453 59 457 62
rect 451 57 457 59
rect 451 55 452 57
rect 454 55 457 57
rect 451 53 457 55
rect 453 42 457 53
rect 461 57 465 59
rect 484 66 488 71
rect 582 73 602 74
rect 582 71 584 73
rect 586 71 602 73
rect 582 70 602 71
rect 484 64 485 66
rect 487 64 488 66
rect 484 62 488 64
rect 493 66 508 67
rect 493 64 495 66
rect 497 65 508 66
rect 497 64 522 65
rect 493 63 518 64
rect 504 62 518 63
rect 520 62 522 64
rect 504 61 522 62
rect 461 55 462 57
rect 464 55 465 57
rect 461 50 465 55
rect 504 50 508 61
rect 501 46 508 50
rect 511 54 515 56
rect 511 52 512 54
rect 514 52 515 54
rect 501 45 505 46
rect 501 43 502 45
rect 504 43 505 45
rect 453 41 493 42
rect 501 41 505 43
rect 511 42 515 52
rect 544 66 562 67
rect 544 64 546 66
rect 548 64 562 66
rect 544 63 562 64
rect 558 57 562 63
rect 558 55 559 57
rect 561 55 562 57
rect 537 50 543 51
rect 453 39 467 41
rect 469 39 493 41
rect 453 38 493 39
rect 509 38 515 42
rect 466 34 470 38
rect 489 34 513 38
rect 558 42 562 55
rect 547 38 562 42
rect 547 34 551 38
rect 565 34 566 45
rect 598 66 602 70
rect 613 67 614 69
rect 598 62 610 66
rect 606 57 610 62
rect 606 55 607 57
rect 609 55 610 57
rect 606 43 610 55
rect 593 40 610 43
rect 593 38 594 40
rect 596 39 610 40
rect 596 38 597 39
rect 335 24 341 33
rect 401 33 407 34
rect 401 31 403 33
rect 405 31 407 33
rect 366 26 372 27
rect 366 24 368 26
rect 370 24 372 26
rect 401 26 407 31
rect 414 32 415 34
rect 417 32 418 34
rect 414 30 418 32
rect 423 33 429 34
rect 423 31 425 33
rect 427 31 429 33
rect 401 24 403 26
rect 405 24 407 26
rect 423 26 429 31
rect 423 24 425 26
rect 427 24 429 26
rect 455 33 461 34
rect 455 31 457 33
rect 459 31 461 33
rect 455 26 461 31
rect 466 32 467 34
rect 469 32 470 34
rect 466 30 470 32
rect 477 33 483 34
rect 477 31 479 33
rect 481 31 483 33
rect 455 24 457 26
rect 459 24 461 26
rect 477 26 483 31
rect 534 33 551 34
rect 534 31 536 33
rect 538 31 551 33
rect 534 30 551 31
rect 582 33 588 34
rect 582 31 584 33
rect 586 31 588 33
rect 477 24 479 26
rect 481 24 483 26
rect 512 26 518 27
rect 512 24 514 26
rect 516 24 518 26
rect 553 26 559 27
rect 553 24 555 26
rect 557 24 559 26
rect 582 24 588 31
rect 593 33 597 38
rect 633 73 637 75
rect 642 74 667 75
rect 751 74 776 75
rect 642 72 644 74
rect 646 73 667 74
rect 646 72 664 73
rect 642 71 664 72
rect 666 71 667 73
rect 643 66 658 67
rect 643 65 654 66
rect 629 64 654 65
rect 656 64 658 66
rect 629 62 631 64
rect 633 63 658 64
rect 663 66 667 71
rect 672 73 682 74
rect 672 71 674 73
rect 676 71 682 73
rect 672 70 682 71
rect 663 64 664 66
rect 666 64 667 66
rect 633 62 647 63
rect 663 62 667 64
rect 629 61 647 62
rect 636 54 640 56
rect 636 52 637 54
rect 639 52 640 54
rect 636 42 640 52
rect 643 50 647 61
rect 678 66 682 70
rect 678 62 698 66
rect 694 59 698 62
rect 686 57 690 59
rect 686 55 687 57
rect 689 55 690 57
rect 686 50 690 55
rect 694 57 700 59
rect 694 55 697 57
rect 699 55 700 57
rect 694 53 700 55
rect 643 46 650 50
rect 646 45 650 46
rect 646 43 647 45
rect 649 43 650 45
rect 636 38 642 42
rect 646 41 650 43
rect 694 42 698 53
rect 658 41 698 42
rect 658 39 682 41
rect 684 39 698 41
rect 658 38 698 39
rect 593 31 594 33
rect 596 31 597 33
rect 593 29 597 31
rect 602 35 608 36
rect 602 33 604 35
rect 606 33 608 35
rect 638 34 662 38
rect 681 34 685 38
rect 736 73 746 74
rect 736 71 742 73
rect 744 71 746 73
rect 736 70 746 71
rect 751 73 772 74
rect 751 71 752 73
rect 754 72 772 73
rect 774 72 776 74
rect 781 73 785 75
rect 754 71 776 72
rect 736 66 740 70
rect 720 62 740 66
rect 720 59 724 62
rect 718 57 724 59
rect 718 55 719 57
rect 721 55 724 57
rect 718 53 724 55
rect 720 42 724 53
rect 728 57 732 59
rect 751 66 755 71
rect 849 73 869 74
rect 849 71 851 73
rect 853 71 869 73
rect 849 70 869 71
rect 751 64 752 66
rect 754 64 755 66
rect 751 62 755 64
rect 760 66 775 67
rect 760 64 762 66
rect 764 65 775 66
rect 764 64 789 65
rect 760 63 785 64
rect 771 62 785 63
rect 787 62 789 64
rect 771 61 789 62
rect 728 55 729 57
rect 731 55 732 57
rect 728 50 732 55
rect 771 50 775 61
rect 768 46 775 50
rect 778 54 782 56
rect 778 52 779 54
rect 781 52 782 54
rect 768 45 772 46
rect 768 43 769 45
rect 771 43 772 45
rect 720 41 760 42
rect 768 41 772 43
rect 778 42 782 52
rect 811 66 829 67
rect 811 64 813 66
rect 815 64 829 66
rect 811 63 829 64
rect 825 57 829 63
rect 825 55 826 57
rect 828 55 829 57
rect 804 50 810 51
rect 720 39 734 41
rect 736 39 760 41
rect 720 38 760 39
rect 776 38 782 42
rect 733 34 737 38
rect 756 34 780 38
rect 825 42 829 55
rect 814 38 829 42
rect 814 34 818 38
rect 832 34 833 45
rect 865 66 869 70
rect 880 67 881 69
rect 865 62 877 66
rect 873 57 877 62
rect 873 55 874 57
rect 876 55 877 57
rect 873 43 877 55
rect 860 40 877 43
rect 860 38 861 40
rect 863 39 877 40
rect 863 38 864 39
rect 602 24 608 33
rect 668 33 674 34
rect 668 31 670 33
rect 672 31 674 33
rect 633 26 639 27
rect 633 24 635 26
rect 637 24 639 26
rect 668 26 674 31
rect 681 32 682 34
rect 684 32 685 34
rect 681 30 685 32
rect 690 33 696 34
rect 690 31 692 33
rect 694 31 696 33
rect 668 24 670 26
rect 672 24 674 26
rect 690 26 696 31
rect 690 24 692 26
rect 694 24 696 26
rect 722 33 728 34
rect 722 31 724 33
rect 726 31 728 33
rect 722 26 728 31
rect 733 32 734 34
rect 736 32 737 34
rect 733 30 737 32
rect 744 33 750 34
rect 744 31 746 33
rect 748 31 750 33
rect 722 24 724 26
rect 726 24 728 26
rect 744 26 750 31
rect 801 33 818 34
rect 801 31 803 33
rect 805 31 818 33
rect 801 30 818 31
rect 849 33 855 34
rect 849 31 851 33
rect 853 31 855 33
rect 744 24 746 26
rect 748 24 750 26
rect 779 26 785 27
rect 779 24 781 26
rect 783 24 785 26
rect 820 26 826 27
rect 820 24 822 26
rect 824 24 826 26
rect 849 24 855 31
rect 860 33 864 38
rect 900 73 904 75
rect 909 74 934 75
rect 1018 74 1043 75
rect 909 72 911 74
rect 913 73 934 74
rect 913 72 931 73
rect 909 71 931 72
rect 933 71 934 73
rect 910 66 925 67
rect 910 65 921 66
rect 896 64 921 65
rect 923 64 925 66
rect 896 62 898 64
rect 900 63 925 64
rect 930 66 934 71
rect 939 73 949 74
rect 939 71 941 73
rect 943 71 949 73
rect 939 70 949 71
rect 930 64 931 66
rect 933 64 934 66
rect 900 62 914 63
rect 930 62 934 64
rect 896 61 914 62
rect 903 54 907 56
rect 903 52 904 54
rect 906 52 907 54
rect 903 42 907 52
rect 910 50 914 61
rect 945 66 949 70
rect 945 62 965 66
rect 961 59 965 62
rect 953 57 957 59
rect 953 55 954 57
rect 956 55 957 57
rect 953 50 957 55
rect 961 57 967 59
rect 961 55 964 57
rect 966 55 967 57
rect 961 53 967 55
rect 910 46 917 50
rect 913 45 917 46
rect 913 43 914 45
rect 916 43 917 45
rect 903 38 909 42
rect 913 41 917 43
rect 961 42 965 53
rect 925 41 965 42
rect 925 39 949 41
rect 951 39 965 41
rect 925 38 965 39
rect 860 31 861 33
rect 863 31 864 33
rect 860 29 864 31
rect 869 35 875 36
rect 869 33 871 35
rect 873 33 875 35
rect 905 34 929 38
rect 948 34 952 38
rect 1003 73 1013 74
rect 1003 71 1009 73
rect 1011 71 1013 73
rect 1003 70 1013 71
rect 1018 73 1039 74
rect 1018 71 1019 73
rect 1021 72 1039 73
rect 1041 72 1043 74
rect 1048 73 1052 75
rect 1021 71 1043 72
rect 1003 66 1007 70
rect 987 62 1007 66
rect 987 59 991 62
rect 985 57 991 59
rect 985 55 986 57
rect 988 55 991 57
rect 985 53 991 55
rect 987 42 991 53
rect 995 57 999 59
rect 1018 66 1022 71
rect 1116 73 1136 74
rect 1116 71 1118 73
rect 1120 71 1136 73
rect 1116 70 1136 71
rect 1018 64 1019 66
rect 1021 64 1022 66
rect 1018 62 1022 64
rect 1027 66 1042 67
rect 1027 64 1029 66
rect 1031 65 1042 66
rect 1031 64 1056 65
rect 1027 63 1052 64
rect 1038 62 1052 63
rect 1054 62 1056 64
rect 1038 61 1056 62
rect 995 55 996 57
rect 998 55 999 57
rect 995 50 999 55
rect 1038 50 1042 61
rect 1035 46 1042 50
rect 1045 54 1049 56
rect 1045 52 1046 54
rect 1048 52 1049 54
rect 1035 45 1039 46
rect 1035 43 1036 45
rect 1038 43 1039 45
rect 987 41 1027 42
rect 1035 41 1039 43
rect 1045 42 1049 52
rect 1078 66 1096 67
rect 1078 64 1080 66
rect 1082 64 1096 66
rect 1078 63 1096 64
rect 1092 57 1096 63
rect 1092 55 1093 57
rect 1095 55 1096 57
rect 1071 50 1077 51
rect 987 39 1001 41
rect 1003 39 1027 41
rect 987 38 1027 39
rect 1043 38 1049 42
rect 1000 34 1004 38
rect 1023 34 1047 38
rect 1092 42 1096 55
rect 1081 38 1096 42
rect 1081 34 1085 38
rect 1099 34 1100 45
rect 1132 66 1136 70
rect 1147 67 1148 69
rect 1132 62 1144 66
rect 1140 57 1144 62
rect 1140 55 1141 57
rect 1143 55 1144 57
rect 1140 43 1144 55
rect 1127 40 1144 43
rect 1127 38 1128 40
rect 1130 39 1144 40
rect 1130 38 1131 39
rect 869 24 875 33
rect 935 33 941 34
rect 935 31 937 33
rect 939 31 941 33
rect 900 26 906 27
rect 900 24 902 26
rect 904 24 906 26
rect 935 26 941 31
rect 948 32 949 34
rect 951 32 952 34
rect 948 30 952 32
rect 957 33 963 34
rect 957 31 959 33
rect 961 31 963 33
rect 935 24 937 26
rect 939 24 941 26
rect 957 26 963 31
rect 957 24 959 26
rect 961 24 963 26
rect 989 33 995 34
rect 989 31 991 33
rect 993 31 995 33
rect 989 26 995 31
rect 1000 32 1001 34
rect 1003 32 1004 34
rect 1000 30 1004 32
rect 1011 33 1017 34
rect 1011 31 1013 33
rect 1015 31 1017 33
rect 989 24 991 26
rect 993 24 995 26
rect 1011 26 1017 31
rect 1068 33 1085 34
rect 1068 31 1070 33
rect 1072 31 1085 33
rect 1068 30 1085 31
rect 1116 33 1122 34
rect 1116 31 1118 33
rect 1120 31 1122 33
rect 1011 24 1013 26
rect 1015 24 1017 26
rect 1046 26 1052 27
rect 1046 24 1048 26
rect 1050 24 1052 26
rect 1087 26 1093 27
rect 1087 24 1089 26
rect 1091 24 1093 26
rect 1116 24 1122 31
rect 1127 33 1131 38
rect 1167 73 1171 75
rect 1176 74 1201 75
rect 1285 74 1310 75
rect 1176 72 1178 74
rect 1180 73 1201 74
rect 1180 72 1198 73
rect 1176 71 1198 72
rect 1200 71 1201 73
rect 1177 66 1192 67
rect 1177 65 1188 66
rect 1163 64 1188 65
rect 1190 64 1192 66
rect 1163 62 1165 64
rect 1167 63 1192 64
rect 1197 66 1201 71
rect 1206 73 1216 74
rect 1206 71 1208 73
rect 1210 71 1216 73
rect 1206 70 1216 71
rect 1197 64 1198 66
rect 1200 64 1201 66
rect 1167 62 1181 63
rect 1197 62 1201 64
rect 1163 61 1181 62
rect 1170 54 1174 56
rect 1170 52 1171 54
rect 1173 52 1174 54
rect 1170 42 1174 52
rect 1177 50 1181 61
rect 1212 66 1216 70
rect 1212 62 1232 66
rect 1228 59 1232 62
rect 1220 57 1224 59
rect 1220 55 1221 57
rect 1223 55 1224 57
rect 1220 50 1224 55
rect 1228 57 1234 59
rect 1228 55 1231 57
rect 1233 55 1234 57
rect 1228 53 1234 55
rect 1177 46 1184 50
rect 1180 45 1184 46
rect 1180 43 1181 45
rect 1183 43 1184 45
rect 1170 38 1176 42
rect 1180 41 1184 43
rect 1228 42 1232 53
rect 1192 41 1232 42
rect 1192 39 1216 41
rect 1218 39 1232 41
rect 1192 38 1232 39
rect 1127 31 1128 33
rect 1130 31 1131 33
rect 1127 29 1131 31
rect 1136 35 1142 36
rect 1136 33 1138 35
rect 1140 33 1142 35
rect 1172 34 1196 38
rect 1215 34 1219 38
rect 1270 73 1280 74
rect 1270 71 1276 73
rect 1278 71 1280 73
rect 1270 70 1280 71
rect 1285 73 1306 74
rect 1285 71 1286 73
rect 1288 72 1306 73
rect 1308 72 1310 74
rect 1315 73 1319 75
rect 1288 71 1310 72
rect 1270 66 1274 70
rect 1254 62 1274 66
rect 1254 59 1258 62
rect 1252 57 1258 59
rect 1252 55 1253 57
rect 1255 55 1258 57
rect 1252 53 1258 55
rect 1254 42 1258 53
rect 1262 57 1266 59
rect 1285 66 1289 71
rect 1383 73 1403 74
rect 1383 71 1385 73
rect 1387 71 1403 73
rect 1383 70 1403 71
rect 1285 64 1286 66
rect 1288 64 1289 66
rect 1285 62 1289 64
rect 1294 66 1309 67
rect 1294 64 1296 66
rect 1298 65 1309 66
rect 1298 64 1323 65
rect 1294 63 1319 64
rect 1305 62 1319 63
rect 1321 62 1323 64
rect 1305 61 1323 62
rect 1262 55 1263 57
rect 1265 55 1266 57
rect 1262 50 1266 55
rect 1305 50 1309 61
rect 1302 46 1309 50
rect 1312 54 1316 56
rect 1312 52 1313 54
rect 1315 52 1316 54
rect 1302 45 1306 46
rect 1302 43 1303 45
rect 1305 43 1306 45
rect 1254 41 1294 42
rect 1302 41 1306 43
rect 1312 42 1316 52
rect 1345 66 1363 67
rect 1345 64 1347 66
rect 1349 64 1363 66
rect 1345 63 1363 64
rect 1359 57 1363 63
rect 1359 55 1360 57
rect 1362 55 1363 57
rect 1338 50 1344 51
rect 1254 39 1268 41
rect 1270 39 1294 41
rect 1254 38 1294 39
rect 1310 38 1316 42
rect 1267 34 1271 38
rect 1290 34 1314 38
rect 1359 42 1363 55
rect 1348 38 1363 42
rect 1348 34 1352 38
rect 1366 34 1367 45
rect 1399 66 1403 70
rect 1414 67 1415 69
rect 1399 62 1411 66
rect 1407 57 1411 62
rect 1407 55 1408 57
rect 1410 55 1411 57
rect 1407 43 1411 55
rect 1394 40 1411 43
rect 1394 38 1395 40
rect 1397 39 1411 40
rect 1397 38 1398 39
rect 1136 24 1142 33
rect 1202 33 1208 34
rect 1202 31 1204 33
rect 1206 31 1208 33
rect 1167 26 1173 27
rect 1167 24 1169 26
rect 1171 24 1173 26
rect 1202 26 1208 31
rect 1215 32 1216 34
rect 1218 32 1219 34
rect 1215 30 1219 32
rect 1224 33 1230 34
rect 1224 31 1226 33
rect 1228 31 1230 33
rect 1202 24 1204 26
rect 1206 24 1208 26
rect 1224 26 1230 31
rect 1224 24 1226 26
rect 1228 24 1230 26
rect 1256 33 1262 34
rect 1256 31 1258 33
rect 1260 31 1262 33
rect 1256 26 1262 31
rect 1267 32 1268 34
rect 1270 32 1271 34
rect 1267 30 1271 32
rect 1278 33 1284 34
rect 1278 31 1280 33
rect 1282 31 1284 33
rect 1256 24 1258 26
rect 1260 24 1262 26
rect 1278 26 1284 31
rect 1335 33 1352 34
rect 1335 31 1337 33
rect 1339 31 1352 33
rect 1335 30 1352 31
rect 1383 33 1389 34
rect 1383 31 1385 33
rect 1387 31 1389 33
rect 1278 24 1280 26
rect 1282 24 1284 26
rect 1313 26 1319 27
rect 1313 24 1315 26
rect 1317 24 1319 26
rect 1354 26 1360 27
rect 1354 24 1356 26
rect 1358 24 1360 26
rect 1383 24 1389 31
rect 1394 33 1398 38
rect 1434 73 1438 75
rect 1443 74 1468 75
rect 1552 74 1577 75
rect 1443 72 1445 74
rect 1447 73 1468 74
rect 1447 72 1465 73
rect 1443 71 1465 72
rect 1467 71 1468 73
rect 1444 66 1459 67
rect 1444 65 1455 66
rect 1430 64 1455 65
rect 1457 64 1459 66
rect 1430 62 1432 64
rect 1434 63 1459 64
rect 1464 66 1468 71
rect 1473 73 1483 74
rect 1473 71 1475 73
rect 1477 71 1483 73
rect 1473 70 1483 71
rect 1464 64 1465 66
rect 1467 64 1468 66
rect 1434 62 1448 63
rect 1464 62 1468 64
rect 1430 61 1448 62
rect 1437 54 1441 56
rect 1437 52 1438 54
rect 1440 52 1441 54
rect 1437 42 1441 52
rect 1444 50 1448 61
rect 1479 66 1483 70
rect 1479 62 1499 66
rect 1495 59 1499 62
rect 1487 57 1491 59
rect 1487 55 1488 57
rect 1490 55 1491 57
rect 1487 50 1491 55
rect 1495 57 1501 59
rect 1495 55 1498 57
rect 1500 55 1501 57
rect 1495 53 1501 55
rect 1444 46 1451 50
rect 1447 45 1451 46
rect 1447 43 1448 45
rect 1450 43 1451 45
rect 1437 38 1443 42
rect 1447 41 1451 43
rect 1495 42 1499 53
rect 1459 41 1499 42
rect 1459 39 1483 41
rect 1485 39 1499 41
rect 1459 38 1499 39
rect 1394 31 1395 33
rect 1397 31 1398 33
rect 1394 29 1398 31
rect 1403 35 1409 36
rect 1403 33 1405 35
rect 1407 33 1409 35
rect 1439 34 1463 38
rect 1482 34 1486 38
rect 1537 73 1547 74
rect 1537 71 1543 73
rect 1545 71 1547 73
rect 1537 70 1547 71
rect 1552 73 1573 74
rect 1552 71 1553 73
rect 1555 72 1573 73
rect 1575 72 1577 74
rect 1582 73 1586 75
rect 1555 71 1577 72
rect 1537 66 1541 70
rect 1521 62 1541 66
rect 1521 59 1525 62
rect 1519 57 1525 59
rect 1519 55 1520 57
rect 1522 55 1525 57
rect 1519 53 1525 55
rect 1521 42 1525 53
rect 1529 57 1533 59
rect 1552 66 1556 71
rect 1650 73 1670 74
rect 1650 71 1652 73
rect 1654 71 1670 73
rect 1650 70 1670 71
rect 1552 64 1553 66
rect 1555 64 1556 66
rect 1552 62 1556 64
rect 1561 66 1576 67
rect 1561 64 1563 66
rect 1565 65 1576 66
rect 1565 64 1590 65
rect 1561 63 1586 64
rect 1572 62 1586 63
rect 1588 62 1590 64
rect 1572 61 1590 62
rect 1529 55 1530 57
rect 1532 55 1533 57
rect 1529 50 1533 55
rect 1572 50 1576 61
rect 1569 46 1576 50
rect 1579 54 1583 56
rect 1579 52 1580 54
rect 1582 52 1583 54
rect 1569 45 1573 46
rect 1569 43 1570 45
rect 1572 43 1573 45
rect 1521 41 1561 42
rect 1569 41 1573 43
rect 1579 42 1583 52
rect 1612 66 1630 67
rect 1612 64 1614 66
rect 1616 64 1630 66
rect 1612 63 1630 64
rect 1626 57 1630 63
rect 1626 55 1627 57
rect 1629 55 1630 57
rect 1605 50 1611 51
rect 1521 39 1535 41
rect 1537 39 1561 41
rect 1521 38 1561 39
rect 1577 38 1583 42
rect 1534 34 1538 38
rect 1557 34 1581 38
rect 1626 42 1630 55
rect 1615 38 1630 42
rect 1615 34 1619 38
rect 1633 34 1634 45
rect 1666 66 1670 70
rect 1681 67 1682 69
rect 1666 62 1678 66
rect 1674 57 1678 62
rect 1674 55 1675 57
rect 1677 55 1678 57
rect 1674 43 1678 55
rect 1661 40 1678 43
rect 1661 38 1662 40
rect 1664 39 1678 40
rect 1664 38 1665 39
rect 1403 24 1409 33
rect 1469 33 1475 34
rect 1469 31 1471 33
rect 1473 31 1475 33
rect 1434 26 1440 27
rect 1434 24 1436 26
rect 1438 24 1440 26
rect 1469 26 1475 31
rect 1482 32 1483 34
rect 1485 32 1486 34
rect 1482 30 1486 32
rect 1491 33 1497 34
rect 1491 31 1493 33
rect 1495 31 1497 33
rect 1469 24 1471 26
rect 1473 24 1475 26
rect 1491 26 1497 31
rect 1491 24 1493 26
rect 1495 24 1497 26
rect 1523 33 1529 34
rect 1523 31 1525 33
rect 1527 31 1529 33
rect 1523 26 1529 31
rect 1534 32 1535 34
rect 1537 32 1538 34
rect 1534 30 1538 32
rect 1545 33 1551 34
rect 1545 31 1547 33
rect 1549 31 1551 33
rect 1523 24 1525 26
rect 1527 24 1529 26
rect 1545 26 1551 31
rect 1602 33 1619 34
rect 1602 31 1604 33
rect 1606 31 1619 33
rect 1602 30 1619 31
rect 1650 33 1656 34
rect 1650 31 1652 33
rect 1654 31 1656 33
rect 1545 24 1547 26
rect 1549 24 1551 26
rect 1580 26 1586 27
rect 1580 24 1582 26
rect 1584 24 1586 26
rect 1621 26 1627 27
rect 1621 24 1623 26
rect 1625 24 1627 26
rect 1650 24 1656 31
rect 1661 33 1665 38
rect 1701 73 1705 75
rect 1710 74 1735 75
rect 1819 74 1844 75
rect 1710 72 1712 74
rect 1714 73 1735 74
rect 1714 72 1732 73
rect 1710 71 1732 72
rect 1734 71 1735 73
rect 1711 66 1726 67
rect 1711 65 1722 66
rect 1697 64 1722 65
rect 1724 64 1726 66
rect 1697 62 1699 64
rect 1701 63 1726 64
rect 1731 66 1735 71
rect 1740 73 1750 74
rect 1740 71 1742 73
rect 1744 71 1750 73
rect 1740 70 1750 71
rect 1731 64 1732 66
rect 1734 64 1735 66
rect 1701 62 1715 63
rect 1731 62 1735 64
rect 1697 61 1715 62
rect 1704 54 1708 56
rect 1704 52 1705 54
rect 1707 52 1708 54
rect 1704 42 1708 52
rect 1711 50 1715 61
rect 1746 66 1750 70
rect 1746 62 1766 66
rect 1762 59 1766 62
rect 1754 57 1758 59
rect 1754 55 1755 57
rect 1757 55 1758 57
rect 1754 50 1758 55
rect 1762 57 1768 59
rect 1762 55 1765 57
rect 1767 55 1768 57
rect 1762 53 1768 55
rect 1711 46 1718 50
rect 1714 45 1718 46
rect 1714 43 1715 45
rect 1717 43 1718 45
rect 1704 38 1710 42
rect 1714 41 1718 43
rect 1762 42 1766 53
rect 1726 41 1766 42
rect 1726 39 1750 41
rect 1752 39 1766 41
rect 1726 38 1766 39
rect 1661 31 1662 33
rect 1664 31 1665 33
rect 1661 29 1665 31
rect 1670 35 1676 36
rect 1670 33 1672 35
rect 1674 33 1676 35
rect 1706 34 1730 38
rect 1749 34 1753 38
rect 1804 73 1814 74
rect 1804 71 1810 73
rect 1812 71 1814 73
rect 1804 70 1814 71
rect 1819 73 1840 74
rect 1819 71 1820 73
rect 1822 72 1840 73
rect 1842 72 1844 74
rect 1849 73 1853 75
rect 1822 71 1844 72
rect 1926 74 1932 80
rect 1987 77 1991 80
rect 2043 78 2045 80
rect 2047 78 2049 80
rect 2043 77 2049 78
rect 2077 78 2079 80
rect 2081 78 2083 80
rect 2077 77 2083 78
rect 2135 77 2139 80
rect 1987 75 1988 77
rect 1990 75 1991 77
rect 2135 75 2136 77
rect 2138 75 2139 77
rect 2155 79 2161 80
rect 2155 77 2157 79
rect 2159 77 2161 79
rect 2155 76 2161 77
rect 2174 79 2180 80
rect 2174 77 2176 79
rect 2178 77 2180 79
rect 2174 76 2180 77
rect 1926 72 1928 74
rect 1930 72 1932 74
rect 1926 71 1932 72
rect 1939 71 1943 73
rect 1804 66 1808 70
rect 1788 62 1808 66
rect 1788 59 1792 62
rect 1786 57 1792 59
rect 1786 55 1787 57
rect 1789 55 1792 57
rect 1786 53 1792 55
rect 1788 42 1792 53
rect 1796 57 1800 59
rect 1819 66 1823 71
rect 1939 69 1940 71
rect 1942 69 1943 71
rect 1819 64 1820 66
rect 1822 64 1823 66
rect 1819 62 1823 64
rect 1828 66 1843 67
rect 1828 64 1830 66
rect 1832 65 1843 66
rect 1832 64 1857 65
rect 1828 63 1853 64
rect 1839 62 1853 63
rect 1855 62 1857 64
rect 1839 61 1857 62
rect 1796 55 1797 57
rect 1799 55 1800 57
rect 1796 50 1800 55
rect 1839 50 1843 61
rect 1836 46 1843 50
rect 1846 54 1850 56
rect 1846 52 1847 54
rect 1849 52 1850 54
rect 1836 45 1840 46
rect 1836 43 1837 45
rect 1839 43 1840 45
rect 1788 41 1828 42
rect 1836 41 1840 43
rect 1846 42 1850 52
rect 1879 66 1897 67
rect 1879 64 1881 66
rect 1883 64 1897 66
rect 1879 63 1897 64
rect 1893 57 1897 63
rect 1893 55 1894 57
rect 1896 55 1897 57
rect 1872 50 1878 51
rect 1788 39 1802 41
rect 1804 39 1828 41
rect 1788 38 1828 39
rect 1844 38 1850 42
rect 1801 34 1805 38
rect 1824 34 1848 38
rect 1893 42 1897 55
rect 1882 38 1897 42
rect 1882 34 1886 38
rect 1900 34 1901 45
rect 1913 66 1917 68
rect 1913 64 1914 66
rect 1916 64 1917 66
rect 1913 58 1917 64
rect 1939 66 1943 69
rect 1939 62 1963 66
rect 1913 54 1924 58
rect 1670 24 1676 33
rect 1736 33 1742 34
rect 1736 31 1738 33
rect 1740 31 1742 33
rect 1701 26 1707 27
rect 1701 24 1703 26
rect 1705 24 1707 26
rect 1736 26 1742 31
rect 1749 32 1750 34
rect 1752 32 1753 34
rect 1749 30 1753 32
rect 1758 33 1764 34
rect 1758 31 1760 33
rect 1762 31 1764 33
rect 1736 24 1738 26
rect 1740 24 1742 26
rect 1758 26 1764 31
rect 1758 24 1760 26
rect 1762 24 1764 26
rect 1790 33 1796 34
rect 1790 31 1792 33
rect 1794 31 1796 33
rect 1790 26 1796 31
rect 1801 32 1802 34
rect 1804 32 1805 34
rect 1801 30 1805 32
rect 1812 33 1818 34
rect 1812 31 1814 33
rect 1816 31 1818 33
rect 1790 24 1792 26
rect 1794 24 1796 26
rect 1812 26 1818 31
rect 1869 33 1886 34
rect 1869 31 1871 33
rect 1873 31 1886 33
rect 1869 30 1886 31
rect 1920 48 1924 54
rect 1959 58 1963 62
rect 1939 57 1955 58
rect 1939 55 1951 57
rect 1953 55 1955 57
rect 1939 54 1955 55
rect 1959 56 1964 58
rect 1959 54 1961 56
rect 1963 54 1964 56
rect 1939 48 1943 54
rect 1959 52 1964 54
rect 1959 50 1963 52
rect 1920 47 1943 48
rect 1920 45 1922 47
rect 1924 45 1943 47
rect 1920 44 1943 45
rect 1931 33 1935 35
rect 1931 31 1932 33
rect 1934 31 1935 33
rect 1812 24 1814 26
rect 1816 24 1818 26
rect 1847 26 1853 27
rect 1847 24 1849 26
rect 1851 24 1853 26
rect 1888 26 1894 27
rect 1888 24 1890 26
rect 1892 24 1894 26
rect 1931 26 1935 31
rect 1939 33 1943 44
rect 1947 47 1963 50
rect 1947 45 1948 47
rect 1950 46 1963 47
rect 1950 45 1951 46
rect 1947 40 1951 45
rect 1947 38 1948 40
rect 1950 38 1951 40
rect 1947 36 1951 38
rect 1987 73 1991 75
rect 1996 74 2021 75
rect 2105 74 2130 75
rect 1996 72 1998 74
rect 2000 73 2021 74
rect 2000 72 2018 73
rect 1996 71 2018 72
rect 2020 71 2021 73
rect 1997 66 2012 67
rect 1997 65 2008 66
rect 1983 64 2008 65
rect 2010 64 2012 66
rect 1983 62 1985 64
rect 1987 63 2012 64
rect 2017 66 2021 71
rect 2026 73 2036 74
rect 2026 71 2028 73
rect 2030 71 2036 73
rect 2026 70 2036 71
rect 2017 64 2018 66
rect 2020 64 2021 66
rect 1987 62 2001 63
rect 2017 62 2021 64
rect 1983 61 2001 62
rect 1990 54 1994 56
rect 1990 52 1991 54
rect 1993 52 1994 54
rect 1990 42 1994 52
rect 1997 50 2001 61
rect 2032 66 2036 70
rect 2032 62 2052 66
rect 2048 59 2052 62
rect 2040 57 2044 59
rect 2040 55 2041 57
rect 2043 55 2044 57
rect 2040 50 2044 55
rect 2048 57 2054 59
rect 2048 55 2051 57
rect 2053 55 2054 57
rect 2048 53 2054 55
rect 1997 46 2004 50
rect 2000 45 2004 46
rect 2000 43 2001 45
rect 2003 43 2004 45
rect 1990 38 1996 42
rect 2000 41 2004 43
rect 2048 42 2052 53
rect 2012 41 2052 42
rect 2012 39 2036 41
rect 2038 39 2052 41
rect 2012 38 2052 39
rect 1992 34 2016 38
rect 2035 34 2039 38
rect 2090 73 2100 74
rect 2090 71 2096 73
rect 2098 71 2100 73
rect 2090 70 2100 71
rect 2105 73 2126 74
rect 2105 71 2106 73
rect 2108 72 2126 73
rect 2128 72 2130 74
rect 2135 73 2139 75
rect 2108 71 2130 72
rect 2199 72 2205 73
rect 2090 66 2094 70
rect 2074 62 2094 66
rect 2074 59 2078 62
rect 2072 57 2078 59
rect 2072 55 2073 57
rect 2075 55 2078 57
rect 2072 53 2078 55
rect 2074 42 2078 53
rect 2082 57 2086 59
rect 2105 66 2109 71
rect 2199 70 2201 72
rect 2203 70 2205 72
rect 2199 69 2205 70
rect 2209 72 2215 80
rect 2209 70 2211 72
rect 2213 70 2215 72
rect 2226 74 2241 75
rect 2226 72 2228 74
rect 2230 72 2241 74
rect 2226 71 2241 72
rect 2209 69 2215 70
rect 2105 64 2106 66
rect 2108 64 2109 66
rect 2105 62 2109 64
rect 2114 66 2129 67
rect 2114 64 2116 66
rect 2118 65 2129 66
rect 2118 64 2143 65
rect 2114 63 2139 64
rect 2125 62 2139 63
rect 2141 62 2143 64
rect 2125 61 2143 62
rect 2082 55 2083 57
rect 2085 55 2086 57
rect 2082 50 2086 55
rect 2125 50 2129 61
rect 2122 46 2129 50
rect 2132 54 2136 56
rect 2132 52 2133 54
rect 2135 52 2136 54
rect 2122 45 2126 46
rect 2122 43 2123 45
rect 2125 43 2126 45
rect 2074 41 2114 42
rect 2122 41 2126 43
rect 2132 42 2136 52
rect 2165 66 2183 67
rect 2165 64 2167 66
rect 2169 64 2183 66
rect 2165 63 2183 64
rect 2179 57 2183 63
rect 2179 55 2180 57
rect 2182 55 2183 57
rect 2158 50 2164 51
rect 2074 39 2088 41
rect 2090 39 2114 41
rect 2074 38 2114 39
rect 2130 38 2136 42
rect 2087 34 2091 38
rect 2110 34 2134 38
rect 2179 42 2183 55
rect 2168 38 2183 42
rect 2168 34 2172 38
rect 2186 34 2187 45
rect 2199 49 2203 69
rect 2237 66 2241 71
rect 2244 74 2248 80
rect 2244 72 2245 74
rect 2247 72 2248 74
rect 2244 70 2248 72
rect 2223 63 2234 65
rect 2223 61 2231 63
rect 2233 61 2234 63
rect 2237 64 2251 66
rect 2237 62 2252 64
rect 2223 59 2234 61
rect 2247 60 2249 62
rect 2251 60 2252 62
rect 2223 49 2227 59
rect 2247 58 2252 60
rect 2199 48 2227 49
rect 2199 46 2201 48
rect 2203 47 2227 48
rect 2203 46 2224 47
rect 2199 45 2224 46
rect 2226 45 2227 47
rect 2243 48 2244 54
rect 2223 43 2227 45
rect 2022 33 2028 34
rect 1939 32 1972 33
rect 1939 30 1968 32
rect 1970 30 1972 32
rect 1939 29 1972 30
rect 2022 31 2024 33
rect 2026 31 2028 33
rect 1931 24 1932 26
rect 1934 24 1935 26
rect 1987 26 1993 27
rect 1987 24 1989 26
rect 1991 24 1993 26
rect 2022 26 2028 31
rect 2035 32 2036 34
rect 2038 32 2039 34
rect 2035 30 2039 32
rect 2044 33 2050 34
rect 2044 31 2046 33
rect 2048 31 2050 33
rect 2022 24 2024 26
rect 2026 24 2028 26
rect 2044 26 2050 31
rect 2044 24 2046 26
rect 2048 24 2050 26
rect 2076 33 2082 34
rect 2076 31 2078 33
rect 2080 31 2082 33
rect 2076 26 2082 31
rect 2087 32 2088 34
rect 2090 32 2091 34
rect 2087 30 2091 32
rect 2098 33 2104 34
rect 2098 31 2100 33
rect 2102 31 2104 33
rect 2076 24 2078 26
rect 2080 24 2082 26
rect 2098 26 2104 31
rect 2155 33 2172 34
rect 2155 31 2157 33
rect 2159 31 2172 33
rect 2155 30 2172 31
rect 2247 41 2251 58
rect 2235 37 2251 41
rect 2226 36 2239 37
rect 2226 34 2228 36
rect 2230 34 2239 36
rect 2267 72 2273 73
rect 2267 70 2269 72
rect 2271 70 2273 72
rect 2267 69 2273 70
rect 2277 72 2283 80
rect 2277 70 2279 72
rect 2281 70 2283 72
rect 2294 74 2309 75
rect 2294 72 2296 74
rect 2298 72 2309 74
rect 2294 71 2309 72
rect 2277 69 2283 70
rect 2267 49 2271 69
rect 2305 66 2309 71
rect 2312 74 2316 80
rect 2312 72 2313 74
rect 2315 72 2316 74
rect 2312 70 2316 72
rect 2291 63 2302 65
rect 2291 61 2299 63
rect 2301 61 2302 63
rect 2305 64 2319 66
rect 2305 62 2320 64
rect 2291 59 2302 61
rect 2315 60 2317 62
rect 2319 60 2320 62
rect 2291 49 2295 59
rect 2315 58 2320 60
rect 2267 48 2295 49
rect 2267 46 2269 48
rect 2271 47 2295 48
rect 2271 46 2292 47
rect 2267 45 2292 46
rect 2294 45 2295 47
rect 2311 48 2312 54
rect 2291 43 2295 45
rect 2226 33 2239 34
rect 2315 41 2319 58
rect 2303 37 2319 41
rect 2294 36 2307 37
rect 2294 34 2296 36
rect 2298 34 2307 36
rect 2294 33 2307 34
rect 2098 24 2100 26
rect 2102 24 2104 26
rect 2133 26 2139 27
rect 2133 24 2135 26
rect 2137 24 2139 26
rect 2174 26 2180 27
rect 2174 24 2176 26
rect 2178 24 2180 26
rect 2210 26 2214 28
rect 2210 24 2211 26
rect 2213 24 2214 26
rect 2243 26 2249 27
rect 2243 24 2245 26
rect 2247 24 2249 26
rect 2278 26 2282 28
rect 2278 24 2279 26
rect 2281 24 2282 26
rect 2311 26 2317 27
rect 2311 24 2313 26
rect 2315 24 2317 26
rect 8 1 14 8
rect 8 -1 10 1
rect 12 -1 14 1
rect 8 -2 14 -1
rect 19 1 23 3
rect 19 -1 20 1
rect 22 -1 23 1
rect 19 -6 23 -1
rect 28 -1 34 8
rect 28 -3 30 -1
rect 32 -3 34 -1
rect 48 1 54 8
rect 48 -1 50 1
rect 52 -1 54 1
rect 48 -2 54 -1
rect 59 1 63 3
rect 59 -1 60 1
rect 62 -1 63 1
rect 28 -4 34 -3
rect 19 -8 20 -6
rect 22 -7 23 -6
rect 22 -8 36 -7
rect 19 -11 36 -8
rect 32 -23 36 -11
rect 32 -25 33 -23
rect 35 -25 36 -23
rect 32 -30 36 -25
rect 24 -34 36 -30
rect 59 -6 63 -1
rect 68 -1 74 8
rect 99 6 101 8
rect 103 6 105 8
rect 99 5 105 6
rect 134 6 136 8
rect 138 6 140 8
rect 68 -3 70 -1
rect 72 -3 74 -1
rect 134 1 140 6
rect 156 6 158 8
rect 160 6 162 8
rect 134 -1 136 1
rect 138 -1 140 1
rect 134 -2 140 -1
rect 147 0 151 2
rect 147 -2 148 0
rect 150 -2 151 0
rect 156 1 162 6
rect 156 -1 158 1
rect 160 -1 162 1
rect 156 -2 162 -1
rect 188 6 190 8
rect 192 6 194 8
rect 188 1 194 6
rect 210 6 212 8
rect 214 6 216 8
rect 188 -1 190 1
rect 192 -1 194 1
rect 188 -2 194 -1
rect 199 0 203 2
rect 199 -2 200 0
rect 202 -2 203 0
rect 210 1 216 6
rect 245 6 247 8
rect 249 6 251 8
rect 245 5 251 6
rect 286 6 288 8
rect 290 6 292 8
rect 286 5 292 6
rect 210 -1 212 1
rect 214 -1 216 1
rect 210 -2 216 -1
rect 267 1 284 2
rect 267 -1 269 1
rect 271 -1 284 1
rect 267 -2 284 -1
rect 315 1 321 8
rect 315 -1 317 1
rect 319 -1 321 1
rect 315 -2 321 -1
rect 326 1 330 3
rect 326 -1 327 1
rect 329 -1 330 1
rect 68 -4 74 -3
rect 59 -8 60 -6
rect 62 -7 63 -6
rect 62 -8 76 -7
rect 59 -11 76 -8
rect 24 -38 28 -34
rect 39 -37 40 -35
rect 72 -23 76 -11
rect 72 -25 73 -23
rect 75 -25 76 -23
rect 72 -30 76 -25
rect 64 -34 76 -30
rect 8 -39 28 -38
rect 8 -41 10 -39
rect 12 -41 28 -39
rect 8 -42 28 -41
rect 64 -38 68 -34
rect 79 -37 80 -35
rect 48 -39 68 -38
rect 48 -41 50 -39
rect 52 -41 68 -39
rect 48 -42 68 -41
rect 104 -6 128 -2
rect 147 -6 151 -2
rect 102 -10 108 -6
rect 124 -7 164 -6
rect 124 -9 148 -7
rect 150 -9 164 -7
rect 102 -20 106 -10
rect 112 -11 116 -9
rect 124 -10 164 -9
rect 112 -13 113 -11
rect 115 -13 116 -11
rect 112 -14 116 -13
rect 102 -22 103 -20
rect 105 -22 106 -20
rect 102 -24 106 -22
rect 109 -18 116 -14
rect 109 -29 113 -18
rect 152 -23 156 -18
rect 152 -25 153 -23
rect 155 -25 156 -23
rect 95 -30 113 -29
rect 95 -32 97 -30
rect 99 -31 113 -30
rect 99 -32 124 -31
rect 95 -33 120 -32
rect 109 -34 120 -33
rect 122 -34 124 -32
rect 109 -35 124 -34
rect 129 -32 133 -30
rect 129 -34 130 -32
rect 132 -34 133 -32
rect 129 -39 133 -34
rect 152 -27 156 -25
rect 160 -21 164 -10
rect 160 -23 166 -21
rect 160 -25 163 -23
rect 165 -25 166 -23
rect 160 -27 166 -25
rect 160 -30 164 -27
rect 144 -34 164 -30
rect 144 -38 148 -34
rect 108 -40 130 -39
rect 99 -43 103 -41
rect 108 -42 110 -40
rect 112 -41 130 -40
rect 132 -41 133 -39
rect 112 -42 133 -41
rect 138 -39 148 -38
rect 138 -41 140 -39
rect 142 -41 148 -39
rect 138 -42 148 -41
rect 199 -6 203 -2
rect 222 -6 246 -2
rect 186 -7 226 -6
rect 186 -9 200 -7
rect 202 -9 226 -7
rect 186 -10 226 -9
rect 186 -21 190 -10
rect 234 -11 238 -9
rect 242 -10 248 -6
rect 234 -13 235 -11
rect 237 -13 238 -11
rect 234 -14 238 -13
rect 234 -18 241 -14
rect 184 -23 190 -21
rect 184 -25 185 -23
rect 187 -25 190 -23
rect 184 -27 190 -25
rect 194 -23 198 -18
rect 194 -25 195 -23
rect 197 -25 198 -23
rect 194 -27 198 -25
rect 186 -30 190 -27
rect 186 -34 206 -30
rect 202 -38 206 -34
rect 237 -29 241 -18
rect 244 -20 248 -10
rect 244 -22 245 -20
rect 247 -22 248 -20
rect 244 -24 248 -22
rect 237 -30 255 -29
rect 217 -32 221 -30
rect 237 -31 251 -30
rect 217 -34 218 -32
rect 220 -34 221 -32
rect 202 -39 212 -38
rect 202 -41 208 -39
rect 210 -41 212 -39
rect 202 -42 212 -41
rect 217 -39 221 -34
rect 226 -32 251 -31
rect 253 -32 255 -30
rect 226 -34 228 -32
rect 230 -33 255 -32
rect 280 -6 284 -2
rect 280 -10 295 -6
rect 270 -19 276 -18
rect 230 -34 241 -33
rect 226 -35 241 -34
rect 291 -23 295 -10
rect 298 -13 299 -2
rect 291 -25 292 -23
rect 294 -25 295 -23
rect 291 -31 295 -25
rect 326 -6 330 -1
rect 335 -1 341 8
rect 366 6 368 8
rect 370 6 372 8
rect 366 5 372 6
rect 401 6 403 8
rect 405 6 407 8
rect 335 -3 337 -1
rect 339 -3 341 -1
rect 401 1 407 6
rect 423 6 425 8
rect 427 6 429 8
rect 401 -1 403 1
rect 405 -1 407 1
rect 401 -2 407 -1
rect 414 0 418 2
rect 414 -2 415 0
rect 417 -2 418 0
rect 423 1 429 6
rect 423 -1 425 1
rect 427 -1 429 1
rect 423 -2 429 -1
rect 455 6 457 8
rect 459 6 461 8
rect 455 1 461 6
rect 477 6 479 8
rect 481 6 483 8
rect 455 -1 457 1
rect 459 -1 461 1
rect 455 -2 461 -1
rect 466 0 470 2
rect 466 -2 467 0
rect 469 -2 470 0
rect 477 1 483 6
rect 512 6 514 8
rect 516 6 518 8
rect 512 5 518 6
rect 553 6 555 8
rect 557 6 559 8
rect 553 5 559 6
rect 477 -1 479 1
rect 481 -1 483 1
rect 477 -2 483 -1
rect 534 1 551 2
rect 534 -1 536 1
rect 538 -1 551 1
rect 534 -2 551 -1
rect 582 1 588 8
rect 582 -1 584 1
rect 586 -1 588 1
rect 582 -2 588 -1
rect 593 1 597 3
rect 593 -1 594 1
rect 596 -1 597 1
rect 335 -4 341 -3
rect 326 -8 327 -6
rect 329 -7 330 -6
rect 329 -8 343 -7
rect 326 -11 343 -8
rect 277 -32 295 -31
rect 277 -34 279 -32
rect 281 -34 295 -32
rect 277 -35 295 -34
rect 339 -23 343 -11
rect 339 -25 340 -23
rect 342 -25 343 -23
rect 339 -30 343 -25
rect 331 -34 343 -30
rect 331 -38 335 -34
rect 346 -37 347 -35
rect 217 -41 218 -39
rect 220 -40 242 -39
rect 220 -41 238 -40
rect 217 -42 238 -41
rect 240 -42 242 -40
rect 108 -43 133 -42
rect 217 -43 242 -42
rect 247 -43 251 -41
rect 315 -39 335 -38
rect 315 -41 317 -39
rect 319 -41 335 -39
rect 315 -42 335 -41
rect 371 -6 395 -2
rect 414 -6 418 -2
rect 369 -10 375 -6
rect 391 -7 431 -6
rect 391 -9 415 -7
rect 417 -9 431 -7
rect 369 -20 373 -10
rect 379 -11 383 -9
rect 391 -10 431 -9
rect 379 -13 380 -11
rect 382 -13 383 -11
rect 379 -14 383 -13
rect 369 -22 370 -20
rect 372 -22 373 -20
rect 369 -24 373 -22
rect 376 -18 383 -14
rect 376 -29 380 -18
rect 419 -23 423 -18
rect 419 -25 420 -23
rect 422 -25 423 -23
rect 362 -30 380 -29
rect 362 -32 364 -30
rect 366 -31 380 -30
rect 366 -32 391 -31
rect 362 -33 387 -32
rect 376 -34 387 -33
rect 389 -34 391 -32
rect 376 -35 391 -34
rect 396 -32 400 -30
rect 396 -34 397 -32
rect 399 -34 400 -32
rect 396 -39 400 -34
rect 419 -27 423 -25
rect 427 -21 431 -10
rect 427 -23 433 -21
rect 427 -25 430 -23
rect 432 -25 433 -23
rect 427 -27 433 -25
rect 427 -30 431 -27
rect 411 -34 431 -30
rect 411 -38 415 -34
rect 375 -40 397 -39
rect 366 -43 370 -41
rect 375 -42 377 -40
rect 379 -41 397 -40
rect 399 -41 400 -39
rect 379 -42 400 -41
rect 405 -39 415 -38
rect 405 -41 407 -39
rect 409 -41 415 -39
rect 405 -42 415 -41
rect 466 -6 470 -2
rect 489 -6 513 -2
rect 453 -7 493 -6
rect 453 -9 467 -7
rect 469 -9 493 -7
rect 453 -10 493 -9
rect 453 -21 457 -10
rect 501 -11 505 -9
rect 509 -10 515 -6
rect 501 -13 502 -11
rect 504 -13 505 -11
rect 501 -14 505 -13
rect 501 -18 508 -14
rect 451 -23 457 -21
rect 451 -25 452 -23
rect 454 -25 457 -23
rect 451 -27 457 -25
rect 461 -23 465 -18
rect 461 -25 462 -23
rect 464 -25 465 -23
rect 461 -27 465 -25
rect 453 -30 457 -27
rect 453 -34 473 -30
rect 469 -38 473 -34
rect 504 -29 508 -18
rect 511 -20 515 -10
rect 511 -22 512 -20
rect 514 -22 515 -20
rect 511 -24 515 -22
rect 504 -30 522 -29
rect 484 -32 488 -30
rect 504 -31 518 -30
rect 484 -34 485 -32
rect 487 -34 488 -32
rect 469 -39 479 -38
rect 469 -41 475 -39
rect 477 -41 479 -39
rect 469 -42 479 -41
rect 484 -39 488 -34
rect 493 -32 518 -31
rect 520 -32 522 -30
rect 493 -34 495 -32
rect 497 -33 522 -32
rect 547 -6 551 -2
rect 547 -10 562 -6
rect 537 -19 543 -18
rect 497 -34 508 -33
rect 493 -35 508 -34
rect 558 -23 562 -10
rect 565 -13 566 -2
rect 558 -25 559 -23
rect 561 -25 562 -23
rect 558 -31 562 -25
rect 593 -6 597 -1
rect 602 -1 608 8
rect 633 6 635 8
rect 637 6 639 8
rect 633 5 639 6
rect 668 6 670 8
rect 672 6 674 8
rect 602 -3 604 -1
rect 606 -3 608 -1
rect 668 1 674 6
rect 690 6 692 8
rect 694 6 696 8
rect 668 -1 670 1
rect 672 -1 674 1
rect 668 -2 674 -1
rect 681 0 685 2
rect 681 -2 682 0
rect 684 -2 685 0
rect 690 1 696 6
rect 690 -1 692 1
rect 694 -1 696 1
rect 690 -2 696 -1
rect 722 6 724 8
rect 726 6 728 8
rect 722 1 728 6
rect 744 6 746 8
rect 748 6 750 8
rect 722 -1 724 1
rect 726 -1 728 1
rect 722 -2 728 -1
rect 733 0 737 2
rect 733 -2 734 0
rect 736 -2 737 0
rect 744 1 750 6
rect 779 6 781 8
rect 783 6 785 8
rect 779 5 785 6
rect 820 6 822 8
rect 824 6 826 8
rect 820 5 826 6
rect 744 -1 746 1
rect 748 -1 750 1
rect 744 -2 750 -1
rect 801 1 818 2
rect 801 -1 803 1
rect 805 -1 818 1
rect 801 -2 818 -1
rect 849 1 855 8
rect 849 -1 851 1
rect 853 -1 855 1
rect 849 -2 855 -1
rect 860 1 864 3
rect 860 -1 861 1
rect 863 -1 864 1
rect 602 -4 608 -3
rect 593 -8 594 -6
rect 596 -7 597 -6
rect 596 -8 610 -7
rect 593 -11 610 -8
rect 544 -32 562 -31
rect 544 -34 546 -32
rect 548 -34 562 -32
rect 544 -35 562 -34
rect 606 -23 610 -11
rect 606 -25 607 -23
rect 609 -25 610 -23
rect 606 -30 610 -25
rect 598 -34 610 -30
rect 598 -38 602 -34
rect 613 -37 614 -35
rect 484 -41 485 -39
rect 487 -40 509 -39
rect 487 -41 505 -40
rect 484 -42 505 -41
rect 507 -42 509 -40
rect 375 -43 400 -42
rect 484 -43 509 -42
rect 514 -43 518 -41
rect 582 -39 602 -38
rect 582 -41 584 -39
rect 586 -41 602 -39
rect 582 -42 602 -41
rect 638 -6 662 -2
rect 681 -6 685 -2
rect 636 -10 642 -6
rect 658 -7 698 -6
rect 658 -9 682 -7
rect 684 -9 698 -7
rect 636 -20 640 -10
rect 646 -11 650 -9
rect 658 -10 698 -9
rect 646 -13 647 -11
rect 649 -13 650 -11
rect 646 -14 650 -13
rect 636 -22 637 -20
rect 639 -22 640 -20
rect 636 -24 640 -22
rect 643 -18 650 -14
rect 643 -29 647 -18
rect 686 -23 690 -18
rect 686 -25 687 -23
rect 689 -25 690 -23
rect 629 -30 647 -29
rect 629 -32 631 -30
rect 633 -31 647 -30
rect 633 -32 658 -31
rect 629 -33 654 -32
rect 643 -34 654 -33
rect 656 -34 658 -32
rect 643 -35 658 -34
rect 663 -32 667 -30
rect 663 -34 664 -32
rect 666 -34 667 -32
rect 663 -39 667 -34
rect 686 -27 690 -25
rect 694 -21 698 -10
rect 694 -23 700 -21
rect 694 -25 697 -23
rect 699 -25 700 -23
rect 694 -27 700 -25
rect 694 -30 698 -27
rect 678 -34 698 -30
rect 678 -38 682 -34
rect 642 -40 664 -39
rect 633 -43 637 -41
rect 642 -42 644 -40
rect 646 -41 664 -40
rect 666 -41 667 -39
rect 646 -42 667 -41
rect 672 -39 682 -38
rect 672 -41 674 -39
rect 676 -41 682 -39
rect 672 -42 682 -41
rect 733 -6 737 -2
rect 756 -6 780 -2
rect 720 -7 760 -6
rect 720 -9 734 -7
rect 736 -9 760 -7
rect 720 -10 760 -9
rect 720 -21 724 -10
rect 768 -11 772 -9
rect 776 -10 782 -6
rect 768 -13 769 -11
rect 771 -13 772 -11
rect 768 -14 772 -13
rect 768 -18 775 -14
rect 718 -23 724 -21
rect 718 -25 719 -23
rect 721 -25 724 -23
rect 718 -27 724 -25
rect 728 -23 732 -18
rect 728 -25 729 -23
rect 731 -25 732 -23
rect 728 -27 732 -25
rect 720 -30 724 -27
rect 720 -34 740 -30
rect 736 -38 740 -34
rect 771 -29 775 -18
rect 778 -20 782 -10
rect 778 -22 779 -20
rect 781 -22 782 -20
rect 778 -24 782 -22
rect 771 -30 789 -29
rect 751 -32 755 -30
rect 771 -31 785 -30
rect 751 -34 752 -32
rect 754 -34 755 -32
rect 736 -39 746 -38
rect 736 -41 742 -39
rect 744 -41 746 -39
rect 736 -42 746 -41
rect 751 -39 755 -34
rect 760 -32 785 -31
rect 787 -32 789 -30
rect 760 -34 762 -32
rect 764 -33 789 -32
rect 814 -6 818 -2
rect 814 -10 829 -6
rect 804 -19 810 -18
rect 764 -34 775 -33
rect 760 -35 775 -34
rect 825 -23 829 -10
rect 832 -13 833 -2
rect 825 -25 826 -23
rect 828 -25 829 -23
rect 825 -31 829 -25
rect 860 -6 864 -1
rect 869 -1 875 8
rect 900 6 902 8
rect 904 6 906 8
rect 900 5 906 6
rect 935 6 937 8
rect 939 6 941 8
rect 869 -3 871 -1
rect 873 -3 875 -1
rect 935 1 941 6
rect 957 6 959 8
rect 961 6 963 8
rect 935 -1 937 1
rect 939 -1 941 1
rect 935 -2 941 -1
rect 948 0 952 2
rect 948 -2 949 0
rect 951 -2 952 0
rect 957 1 963 6
rect 957 -1 959 1
rect 961 -1 963 1
rect 957 -2 963 -1
rect 989 6 991 8
rect 993 6 995 8
rect 989 1 995 6
rect 1011 6 1013 8
rect 1015 6 1017 8
rect 989 -1 991 1
rect 993 -1 995 1
rect 989 -2 995 -1
rect 1000 0 1004 2
rect 1000 -2 1001 0
rect 1003 -2 1004 0
rect 1011 1 1017 6
rect 1046 6 1048 8
rect 1050 6 1052 8
rect 1046 5 1052 6
rect 1087 6 1089 8
rect 1091 6 1093 8
rect 1087 5 1093 6
rect 1011 -1 1013 1
rect 1015 -1 1017 1
rect 1011 -2 1017 -1
rect 1068 1 1085 2
rect 1068 -1 1070 1
rect 1072 -1 1085 1
rect 1068 -2 1085 -1
rect 1116 1 1122 8
rect 1116 -1 1118 1
rect 1120 -1 1122 1
rect 1116 -2 1122 -1
rect 1127 1 1131 3
rect 1127 -1 1128 1
rect 1130 -1 1131 1
rect 869 -4 875 -3
rect 860 -8 861 -6
rect 863 -7 864 -6
rect 863 -8 877 -7
rect 860 -11 877 -8
rect 811 -32 829 -31
rect 811 -34 813 -32
rect 815 -34 829 -32
rect 811 -35 829 -34
rect 873 -23 877 -11
rect 873 -25 874 -23
rect 876 -25 877 -23
rect 873 -30 877 -25
rect 865 -34 877 -30
rect 865 -38 869 -34
rect 880 -37 881 -35
rect 751 -41 752 -39
rect 754 -40 776 -39
rect 754 -41 772 -40
rect 751 -42 772 -41
rect 774 -42 776 -40
rect 642 -43 667 -42
rect 751 -43 776 -42
rect 781 -43 785 -41
rect 849 -39 869 -38
rect 849 -41 851 -39
rect 853 -41 869 -39
rect 849 -42 869 -41
rect 905 -6 929 -2
rect 948 -6 952 -2
rect 903 -10 909 -6
rect 925 -7 965 -6
rect 925 -9 949 -7
rect 951 -9 965 -7
rect 903 -20 907 -10
rect 913 -11 917 -9
rect 925 -10 965 -9
rect 913 -13 914 -11
rect 916 -13 917 -11
rect 913 -14 917 -13
rect 903 -22 904 -20
rect 906 -22 907 -20
rect 903 -24 907 -22
rect 910 -18 917 -14
rect 910 -29 914 -18
rect 953 -23 957 -18
rect 953 -25 954 -23
rect 956 -25 957 -23
rect 896 -30 914 -29
rect 896 -32 898 -30
rect 900 -31 914 -30
rect 900 -32 925 -31
rect 896 -33 921 -32
rect 910 -34 921 -33
rect 923 -34 925 -32
rect 910 -35 925 -34
rect 930 -32 934 -30
rect 930 -34 931 -32
rect 933 -34 934 -32
rect 930 -39 934 -34
rect 953 -27 957 -25
rect 961 -21 965 -10
rect 961 -23 967 -21
rect 961 -25 964 -23
rect 966 -25 967 -23
rect 961 -27 967 -25
rect 961 -30 965 -27
rect 945 -34 965 -30
rect 945 -38 949 -34
rect 909 -40 931 -39
rect 900 -43 904 -41
rect 909 -42 911 -40
rect 913 -41 931 -40
rect 933 -41 934 -39
rect 913 -42 934 -41
rect 939 -39 949 -38
rect 939 -41 941 -39
rect 943 -41 949 -39
rect 939 -42 949 -41
rect 1000 -6 1004 -2
rect 1023 -6 1047 -2
rect 987 -7 1027 -6
rect 987 -9 1001 -7
rect 1003 -9 1027 -7
rect 987 -10 1027 -9
rect 987 -21 991 -10
rect 1035 -11 1039 -9
rect 1043 -10 1049 -6
rect 1035 -13 1036 -11
rect 1038 -13 1039 -11
rect 1035 -14 1039 -13
rect 1035 -18 1042 -14
rect 985 -23 991 -21
rect 985 -25 986 -23
rect 988 -25 991 -23
rect 985 -27 991 -25
rect 995 -23 999 -18
rect 995 -25 996 -23
rect 998 -25 999 -23
rect 995 -27 999 -25
rect 987 -30 991 -27
rect 987 -34 1007 -30
rect 1003 -38 1007 -34
rect 1038 -29 1042 -18
rect 1045 -20 1049 -10
rect 1045 -22 1046 -20
rect 1048 -22 1049 -20
rect 1045 -24 1049 -22
rect 1038 -30 1056 -29
rect 1018 -32 1022 -30
rect 1038 -31 1052 -30
rect 1018 -34 1019 -32
rect 1021 -34 1022 -32
rect 1003 -39 1013 -38
rect 1003 -41 1009 -39
rect 1011 -41 1013 -39
rect 1003 -42 1013 -41
rect 1018 -39 1022 -34
rect 1027 -32 1052 -31
rect 1054 -32 1056 -30
rect 1027 -34 1029 -32
rect 1031 -33 1056 -32
rect 1081 -6 1085 -2
rect 1081 -10 1096 -6
rect 1071 -19 1077 -18
rect 1031 -34 1042 -33
rect 1027 -35 1042 -34
rect 1092 -23 1096 -10
rect 1099 -13 1100 -2
rect 1092 -25 1093 -23
rect 1095 -25 1096 -23
rect 1092 -31 1096 -25
rect 1127 -6 1131 -1
rect 1136 -1 1142 8
rect 1167 6 1169 8
rect 1171 6 1173 8
rect 1167 5 1173 6
rect 1202 6 1204 8
rect 1206 6 1208 8
rect 1136 -3 1138 -1
rect 1140 -3 1142 -1
rect 1202 1 1208 6
rect 1224 6 1226 8
rect 1228 6 1230 8
rect 1202 -1 1204 1
rect 1206 -1 1208 1
rect 1202 -2 1208 -1
rect 1215 0 1219 2
rect 1215 -2 1216 0
rect 1218 -2 1219 0
rect 1224 1 1230 6
rect 1224 -1 1226 1
rect 1228 -1 1230 1
rect 1224 -2 1230 -1
rect 1256 6 1258 8
rect 1260 6 1262 8
rect 1256 1 1262 6
rect 1278 6 1280 8
rect 1282 6 1284 8
rect 1256 -1 1258 1
rect 1260 -1 1262 1
rect 1256 -2 1262 -1
rect 1267 0 1271 2
rect 1267 -2 1268 0
rect 1270 -2 1271 0
rect 1278 1 1284 6
rect 1313 6 1315 8
rect 1317 6 1319 8
rect 1313 5 1319 6
rect 1354 6 1356 8
rect 1358 6 1360 8
rect 1354 5 1360 6
rect 1278 -1 1280 1
rect 1282 -1 1284 1
rect 1278 -2 1284 -1
rect 1335 1 1352 2
rect 1335 -1 1337 1
rect 1339 -1 1352 1
rect 1335 -2 1352 -1
rect 1383 1 1389 8
rect 1383 -1 1385 1
rect 1387 -1 1389 1
rect 1383 -2 1389 -1
rect 1394 1 1398 3
rect 1394 -1 1395 1
rect 1397 -1 1398 1
rect 1136 -4 1142 -3
rect 1127 -8 1128 -6
rect 1130 -7 1131 -6
rect 1130 -8 1144 -7
rect 1127 -11 1144 -8
rect 1078 -32 1096 -31
rect 1078 -34 1080 -32
rect 1082 -34 1096 -32
rect 1078 -35 1096 -34
rect 1140 -23 1144 -11
rect 1140 -25 1141 -23
rect 1143 -25 1144 -23
rect 1140 -30 1144 -25
rect 1132 -34 1144 -30
rect 1132 -38 1136 -34
rect 1147 -37 1148 -35
rect 1018 -41 1019 -39
rect 1021 -40 1043 -39
rect 1021 -41 1039 -40
rect 1018 -42 1039 -41
rect 1041 -42 1043 -40
rect 909 -43 934 -42
rect 1018 -43 1043 -42
rect 1048 -43 1052 -41
rect 1116 -39 1136 -38
rect 1116 -41 1118 -39
rect 1120 -41 1136 -39
rect 1116 -42 1136 -41
rect 1172 -6 1196 -2
rect 1215 -6 1219 -2
rect 1170 -10 1176 -6
rect 1192 -7 1232 -6
rect 1192 -9 1216 -7
rect 1218 -9 1232 -7
rect 1170 -20 1174 -10
rect 1180 -11 1184 -9
rect 1192 -10 1232 -9
rect 1180 -13 1181 -11
rect 1183 -13 1184 -11
rect 1180 -14 1184 -13
rect 1170 -22 1171 -20
rect 1173 -22 1174 -20
rect 1170 -24 1174 -22
rect 1177 -18 1184 -14
rect 1177 -29 1181 -18
rect 1220 -23 1224 -18
rect 1220 -25 1221 -23
rect 1223 -25 1224 -23
rect 1163 -30 1181 -29
rect 1163 -32 1165 -30
rect 1167 -31 1181 -30
rect 1167 -32 1192 -31
rect 1163 -33 1188 -32
rect 1177 -34 1188 -33
rect 1190 -34 1192 -32
rect 1177 -35 1192 -34
rect 1197 -32 1201 -30
rect 1197 -34 1198 -32
rect 1200 -34 1201 -32
rect 1197 -39 1201 -34
rect 1220 -27 1224 -25
rect 1228 -21 1232 -10
rect 1228 -23 1234 -21
rect 1228 -25 1231 -23
rect 1233 -25 1234 -23
rect 1228 -27 1234 -25
rect 1228 -30 1232 -27
rect 1212 -34 1232 -30
rect 1212 -38 1216 -34
rect 1176 -40 1198 -39
rect 1167 -43 1171 -41
rect 1176 -42 1178 -40
rect 1180 -41 1198 -40
rect 1200 -41 1201 -39
rect 1180 -42 1201 -41
rect 1206 -39 1216 -38
rect 1206 -41 1208 -39
rect 1210 -41 1216 -39
rect 1206 -42 1216 -41
rect 1267 -6 1271 -2
rect 1290 -6 1314 -2
rect 1254 -7 1294 -6
rect 1254 -9 1268 -7
rect 1270 -9 1294 -7
rect 1254 -10 1294 -9
rect 1254 -21 1258 -10
rect 1302 -11 1306 -9
rect 1310 -10 1316 -6
rect 1302 -13 1303 -11
rect 1305 -13 1306 -11
rect 1302 -14 1306 -13
rect 1302 -18 1309 -14
rect 1252 -23 1258 -21
rect 1252 -25 1253 -23
rect 1255 -25 1258 -23
rect 1252 -27 1258 -25
rect 1262 -23 1266 -18
rect 1262 -25 1263 -23
rect 1265 -25 1266 -23
rect 1262 -27 1266 -25
rect 1254 -30 1258 -27
rect 1254 -34 1274 -30
rect 1270 -38 1274 -34
rect 1305 -29 1309 -18
rect 1312 -20 1316 -10
rect 1312 -22 1313 -20
rect 1315 -22 1316 -20
rect 1312 -24 1316 -22
rect 1305 -30 1323 -29
rect 1285 -32 1289 -30
rect 1305 -31 1319 -30
rect 1285 -34 1286 -32
rect 1288 -34 1289 -32
rect 1270 -39 1280 -38
rect 1270 -41 1276 -39
rect 1278 -41 1280 -39
rect 1270 -42 1280 -41
rect 1285 -39 1289 -34
rect 1294 -32 1319 -31
rect 1321 -32 1323 -30
rect 1294 -34 1296 -32
rect 1298 -33 1323 -32
rect 1348 -6 1352 -2
rect 1348 -10 1363 -6
rect 1338 -19 1344 -18
rect 1298 -34 1309 -33
rect 1294 -35 1309 -34
rect 1359 -23 1363 -10
rect 1366 -13 1367 -2
rect 1359 -25 1360 -23
rect 1362 -25 1363 -23
rect 1359 -31 1363 -25
rect 1394 -6 1398 -1
rect 1403 -1 1409 8
rect 1434 6 1436 8
rect 1438 6 1440 8
rect 1434 5 1440 6
rect 1469 6 1471 8
rect 1473 6 1475 8
rect 1403 -3 1405 -1
rect 1407 -3 1409 -1
rect 1469 1 1475 6
rect 1491 6 1493 8
rect 1495 6 1497 8
rect 1469 -1 1471 1
rect 1473 -1 1475 1
rect 1469 -2 1475 -1
rect 1482 0 1486 2
rect 1482 -2 1483 0
rect 1485 -2 1486 0
rect 1491 1 1497 6
rect 1491 -1 1493 1
rect 1495 -1 1497 1
rect 1491 -2 1497 -1
rect 1523 6 1525 8
rect 1527 6 1529 8
rect 1523 1 1529 6
rect 1545 6 1547 8
rect 1549 6 1551 8
rect 1523 -1 1525 1
rect 1527 -1 1529 1
rect 1523 -2 1529 -1
rect 1534 0 1538 2
rect 1534 -2 1535 0
rect 1537 -2 1538 0
rect 1545 1 1551 6
rect 1580 6 1582 8
rect 1584 6 1586 8
rect 1580 5 1586 6
rect 1621 6 1623 8
rect 1625 6 1627 8
rect 1621 5 1627 6
rect 1545 -1 1547 1
rect 1549 -1 1551 1
rect 1545 -2 1551 -1
rect 1602 1 1619 2
rect 1602 -1 1604 1
rect 1606 -1 1619 1
rect 1602 -2 1619 -1
rect 1650 1 1656 8
rect 1650 -1 1652 1
rect 1654 -1 1656 1
rect 1650 -2 1656 -1
rect 1661 1 1665 3
rect 1661 -1 1662 1
rect 1664 -1 1665 1
rect 1403 -4 1409 -3
rect 1394 -8 1395 -6
rect 1397 -7 1398 -6
rect 1397 -8 1411 -7
rect 1394 -11 1411 -8
rect 1345 -32 1363 -31
rect 1345 -34 1347 -32
rect 1349 -34 1363 -32
rect 1345 -35 1363 -34
rect 1407 -23 1411 -11
rect 1407 -25 1408 -23
rect 1410 -25 1411 -23
rect 1407 -30 1411 -25
rect 1399 -34 1411 -30
rect 1399 -38 1403 -34
rect 1414 -37 1415 -35
rect 1285 -41 1286 -39
rect 1288 -40 1310 -39
rect 1288 -41 1306 -40
rect 1285 -42 1306 -41
rect 1308 -42 1310 -40
rect 1176 -43 1201 -42
rect 1285 -43 1310 -42
rect 1315 -43 1319 -41
rect 1383 -39 1403 -38
rect 1383 -41 1385 -39
rect 1387 -41 1403 -39
rect 1383 -42 1403 -41
rect 1439 -6 1463 -2
rect 1482 -6 1486 -2
rect 1437 -10 1443 -6
rect 1459 -7 1499 -6
rect 1459 -9 1483 -7
rect 1485 -9 1499 -7
rect 1437 -20 1441 -10
rect 1447 -11 1451 -9
rect 1459 -10 1499 -9
rect 1447 -13 1448 -11
rect 1450 -13 1451 -11
rect 1447 -14 1451 -13
rect 1437 -22 1438 -20
rect 1440 -22 1441 -20
rect 1437 -24 1441 -22
rect 1444 -18 1451 -14
rect 1444 -29 1448 -18
rect 1487 -23 1491 -18
rect 1487 -25 1488 -23
rect 1490 -25 1491 -23
rect 1430 -30 1448 -29
rect 1430 -32 1432 -30
rect 1434 -31 1448 -30
rect 1434 -32 1459 -31
rect 1430 -33 1455 -32
rect 1444 -34 1455 -33
rect 1457 -34 1459 -32
rect 1444 -35 1459 -34
rect 1464 -32 1468 -30
rect 1464 -34 1465 -32
rect 1467 -34 1468 -32
rect 1464 -39 1468 -34
rect 1487 -27 1491 -25
rect 1495 -21 1499 -10
rect 1495 -23 1501 -21
rect 1495 -25 1498 -23
rect 1500 -25 1501 -23
rect 1495 -27 1501 -25
rect 1495 -30 1499 -27
rect 1479 -34 1499 -30
rect 1479 -38 1483 -34
rect 1443 -40 1465 -39
rect 1434 -43 1438 -41
rect 1443 -42 1445 -40
rect 1447 -41 1465 -40
rect 1467 -41 1468 -39
rect 1447 -42 1468 -41
rect 1473 -39 1483 -38
rect 1473 -41 1475 -39
rect 1477 -41 1483 -39
rect 1473 -42 1483 -41
rect 1534 -6 1538 -2
rect 1557 -6 1581 -2
rect 1521 -7 1561 -6
rect 1521 -9 1535 -7
rect 1537 -9 1561 -7
rect 1521 -10 1561 -9
rect 1521 -21 1525 -10
rect 1569 -11 1573 -9
rect 1577 -10 1583 -6
rect 1569 -13 1570 -11
rect 1572 -13 1573 -11
rect 1569 -14 1573 -13
rect 1569 -18 1576 -14
rect 1519 -23 1525 -21
rect 1519 -25 1520 -23
rect 1522 -25 1525 -23
rect 1519 -27 1525 -25
rect 1529 -23 1533 -18
rect 1529 -25 1530 -23
rect 1532 -25 1533 -23
rect 1529 -27 1533 -25
rect 1521 -30 1525 -27
rect 1521 -34 1541 -30
rect 1537 -38 1541 -34
rect 1572 -29 1576 -18
rect 1579 -20 1583 -10
rect 1579 -22 1580 -20
rect 1582 -22 1583 -20
rect 1579 -24 1583 -22
rect 1572 -30 1590 -29
rect 1552 -32 1556 -30
rect 1572 -31 1586 -30
rect 1552 -34 1553 -32
rect 1555 -34 1556 -32
rect 1537 -39 1547 -38
rect 1537 -41 1543 -39
rect 1545 -41 1547 -39
rect 1537 -42 1547 -41
rect 1552 -39 1556 -34
rect 1561 -32 1586 -31
rect 1588 -32 1590 -30
rect 1561 -34 1563 -32
rect 1565 -33 1590 -32
rect 1615 -6 1619 -2
rect 1615 -10 1630 -6
rect 1605 -19 1611 -18
rect 1565 -34 1576 -33
rect 1561 -35 1576 -34
rect 1626 -23 1630 -10
rect 1633 -13 1634 -2
rect 1626 -25 1627 -23
rect 1629 -25 1630 -23
rect 1626 -31 1630 -25
rect 1661 -6 1665 -1
rect 1670 -1 1676 8
rect 1701 6 1703 8
rect 1705 6 1707 8
rect 1701 5 1707 6
rect 1736 6 1738 8
rect 1740 6 1742 8
rect 1670 -3 1672 -1
rect 1674 -3 1676 -1
rect 1736 1 1742 6
rect 1758 6 1760 8
rect 1762 6 1764 8
rect 1736 -1 1738 1
rect 1740 -1 1742 1
rect 1736 -2 1742 -1
rect 1749 0 1753 2
rect 1749 -2 1750 0
rect 1752 -2 1753 0
rect 1758 1 1764 6
rect 1758 -1 1760 1
rect 1762 -1 1764 1
rect 1758 -2 1764 -1
rect 1790 6 1792 8
rect 1794 6 1796 8
rect 1790 1 1796 6
rect 1812 6 1814 8
rect 1816 6 1818 8
rect 1790 -1 1792 1
rect 1794 -1 1796 1
rect 1790 -2 1796 -1
rect 1801 0 1805 2
rect 1801 -2 1802 0
rect 1804 -2 1805 0
rect 1812 1 1818 6
rect 1847 6 1849 8
rect 1851 6 1853 8
rect 1847 5 1853 6
rect 1888 6 1890 8
rect 1892 6 1894 8
rect 1888 5 1894 6
rect 1931 6 1932 8
rect 1934 6 1935 8
rect 1812 -1 1814 1
rect 1816 -1 1818 1
rect 1812 -2 1818 -1
rect 1869 1 1886 2
rect 1869 -1 1871 1
rect 1873 -1 1886 1
rect 1869 -2 1886 -1
rect 1670 -4 1676 -3
rect 1661 -8 1662 -6
rect 1664 -7 1665 -6
rect 1664 -8 1678 -7
rect 1661 -11 1678 -8
rect 1612 -32 1630 -31
rect 1612 -34 1614 -32
rect 1616 -34 1630 -32
rect 1612 -35 1630 -34
rect 1674 -23 1678 -11
rect 1674 -25 1675 -23
rect 1677 -25 1678 -23
rect 1674 -30 1678 -25
rect 1666 -34 1678 -30
rect 1666 -38 1670 -34
rect 1681 -37 1682 -35
rect 1552 -41 1553 -39
rect 1555 -40 1577 -39
rect 1555 -41 1573 -40
rect 1552 -42 1573 -41
rect 1575 -42 1577 -40
rect 1443 -43 1468 -42
rect 1552 -43 1577 -42
rect 1582 -43 1586 -41
rect 1650 -39 1670 -38
rect 1650 -41 1652 -39
rect 1654 -41 1670 -39
rect 1650 -42 1670 -41
rect 1706 -6 1730 -2
rect 1749 -6 1753 -2
rect 1704 -10 1710 -6
rect 1726 -7 1766 -6
rect 1726 -9 1750 -7
rect 1752 -9 1766 -7
rect 1704 -20 1708 -10
rect 1714 -11 1718 -9
rect 1726 -10 1766 -9
rect 1714 -13 1715 -11
rect 1717 -13 1718 -11
rect 1714 -14 1718 -13
rect 1704 -22 1705 -20
rect 1707 -22 1708 -20
rect 1704 -24 1708 -22
rect 1711 -18 1718 -14
rect 1711 -29 1715 -18
rect 1754 -23 1758 -18
rect 1754 -25 1755 -23
rect 1757 -25 1758 -23
rect 1697 -30 1715 -29
rect 1697 -32 1699 -30
rect 1701 -31 1715 -30
rect 1701 -32 1726 -31
rect 1697 -33 1722 -32
rect 1711 -34 1722 -33
rect 1724 -34 1726 -32
rect 1711 -35 1726 -34
rect 1731 -32 1735 -30
rect 1731 -34 1732 -32
rect 1734 -34 1735 -32
rect 1731 -39 1735 -34
rect 1754 -27 1758 -25
rect 1762 -21 1766 -10
rect 1762 -23 1768 -21
rect 1762 -25 1765 -23
rect 1767 -25 1768 -23
rect 1762 -27 1768 -25
rect 1762 -30 1766 -27
rect 1746 -34 1766 -30
rect 1746 -38 1750 -34
rect 1710 -40 1732 -39
rect 1701 -43 1705 -41
rect 1710 -42 1712 -40
rect 1714 -41 1732 -40
rect 1734 -41 1735 -39
rect 1714 -42 1735 -41
rect 1740 -39 1750 -38
rect 1740 -41 1742 -39
rect 1744 -41 1750 -39
rect 1740 -42 1750 -41
rect 1801 -6 1805 -2
rect 1824 -6 1848 -2
rect 1788 -7 1828 -6
rect 1788 -9 1802 -7
rect 1804 -9 1828 -7
rect 1788 -10 1828 -9
rect 1788 -21 1792 -10
rect 1836 -11 1840 -9
rect 1844 -10 1850 -6
rect 1836 -13 1837 -11
rect 1839 -13 1840 -11
rect 1836 -14 1840 -13
rect 1836 -18 1843 -14
rect 1786 -23 1792 -21
rect 1786 -25 1787 -23
rect 1789 -25 1792 -23
rect 1786 -27 1792 -25
rect 1796 -23 1800 -18
rect 1796 -25 1797 -23
rect 1799 -25 1800 -23
rect 1796 -27 1800 -25
rect 1788 -30 1792 -27
rect 1788 -34 1808 -30
rect 1804 -38 1808 -34
rect 1839 -29 1843 -18
rect 1846 -20 1850 -10
rect 1846 -22 1847 -20
rect 1849 -22 1850 -20
rect 1846 -24 1850 -22
rect 1839 -30 1857 -29
rect 1819 -32 1823 -30
rect 1839 -31 1853 -30
rect 1819 -34 1820 -32
rect 1822 -34 1823 -32
rect 1804 -39 1814 -38
rect 1804 -41 1810 -39
rect 1812 -41 1814 -39
rect 1804 -42 1814 -41
rect 1819 -39 1823 -34
rect 1828 -32 1853 -31
rect 1855 -32 1857 -30
rect 1828 -34 1830 -32
rect 1832 -33 1857 -32
rect 1882 -6 1886 -2
rect 1882 -10 1897 -6
rect 1872 -19 1878 -18
rect 1832 -34 1843 -33
rect 1828 -35 1843 -34
rect 1893 -23 1897 -10
rect 1900 -13 1901 -2
rect 1893 -25 1894 -23
rect 1896 -25 1897 -23
rect 1893 -31 1897 -25
rect 1931 1 1935 6
rect 1987 6 1989 8
rect 1991 6 1993 8
rect 1987 5 1993 6
rect 2022 6 2024 8
rect 2026 6 2028 8
rect 1931 -1 1932 1
rect 1934 -1 1935 1
rect 1931 -3 1935 -1
rect 1939 2 1972 3
rect 1939 0 1968 2
rect 1970 0 1972 2
rect 1939 -1 1972 0
rect 2022 1 2028 6
rect 2044 6 2046 8
rect 2048 6 2050 8
rect 2022 -1 2024 1
rect 2026 -1 2028 1
rect 1939 -12 1943 -1
rect 2022 -2 2028 -1
rect 2035 0 2039 2
rect 2035 -2 2036 0
rect 2038 -2 2039 0
rect 2044 1 2050 6
rect 2044 -1 2046 1
rect 2048 -1 2050 1
rect 2044 -2 2050 -1
rect 2076 6 2078 8
rect 2080 6 2082 8
rect 2076 1 2082 6
rect 2098 6 2100 8
rect 2102 6 2104 8
rect 2076 -1 2078 1
rect 2080 -1 2082 1
rect 2076 -2 2082 -1
rect 2087 0 2091 2
rect 2087 -2 2088 0
rect 2090 -2 2091 0
rect 2098 1 2104 6
rect 2133 6 2135 8
rect 2137 6 2139 8
rect 2133 5 2139 6
rect 2174 6 2176 8
rect 2178 6 2180 8
rect 2174 5 2180 6
rect 2210 6 2211 8
rect 2213 6 2214 8
rect 2210 4 2214 6
rect 2243 6 2245 8
rect 2247 6 2249 8
rect 2243 5 2249 6
rect 2278 6 2279 8
rect 2281 6 2282 8
rect 2278 4 2282 6
rect 2311 6 2313 8
rect 2315 6 2317 8
rect 2311 5 2317 6
rect 2098 -1 2100 1
rect 2102 -1 2104 1
rect 2098 -2 2104 -1
rect 2155 1 2172 2
rect 2155 -1 2157 1
rect 2159 -1 2172 1
rect 2155 -2 2172 -1
rect 1920 -13 1943 -12
rect 1920 -15 1922 -13
rect 1924 -15 1943 -13
rect 1920 -16 1943 -15
rect 1920 -22 1924 -16
rect 1879 -32 1897 -31
rect 1879 -34 1881 -32
rect 1883 -34 1897 -32
rect 1879 -35 1897 -34
rect 1913 -26 1924 -22
rect 1913 -32 1917 -26
rect 1939 -22 1943 -16
rect 1947 -6 1951 -4
rect 1947 -8 1948 -6
rect 1950 -8 1951 -6
rect 1947 -13 1951 -8
rect 1947 -15 1948 -13
rect 1950 -14 1951 -13
rect 1950 -15 1963 -14
rect 1947 -18 1963 -15
rect 1959 -20 1963 -18
rect 1959 -22 1964 -20
rect 1939 -23 1955 -22
rect 1939 -25 1951 -23
rect 1953 -25 1955 -23
rect 1939 -26 1955 -25
rect 1959 -24 1961 -22
rect 1963 -24 1964 -22
rect 1959 -26 1964 -24
rect 1913 -34 1914 -32
rect 1916 -34 1917 -32
rect 1913 -36 1917 -34
rect 1959 -30 1963 -26
rect 1939 -34 1963 -30
rect 1939 -37 1943 -34
rect 1939 -39 1940 -37
rect 1942 -39 1943 -37
rect 1819 -41 1820 -39
rect 1822 -40 1844 -39
rect 1822 -41 1840 -40
rect 1819 -42 1840 -41
rect 1842 -42 1844 -40
rect 1710 -43 1735 -42
rect 1819 -43 1844 -42
rect 1849 -43 1853 -41
rect 1926 -40 1932 -39
rect 1926 -42 1928 -40
rect 1930 -42 1932 -40
rect 1939 -41 1943 -39
rect 1992 -6 2016 -2
rect 2035 -6 2039 -2
rect 1990 -10 1996 -6
rect 2012 -7 2052 -6
rect 2012 -9 2036 -7
rect 2038 -9 2052 -7
rect 1990 -20 1994 -10
rect 2000 -11 2004 -9
rect 2012 -10 2052 -9
rect 2000 -13 2001 -11
rect 2003 -13 2004 -11
rect 2000 -14 2004 -13
rect 1990 -22 1991 -20
rect 1993 -22 1994 -20
rect 1990 -24 1994 -22
rect 1997 -18 2004 -14
rect 1997 -29 2001 -18
rect 2040 -23 2044 -18
rect 2040 -25 2041 -23
rect 2043 -25 2044 -23
rect 1983 -30 2001 -29
rect 1983 -32 1985 -30
rect 1987 -31 2001 -30
rect 1987 -32 2012 -31
rect 1983 -33 2008 -32
rect 1997 -34 2008 -33
rect 2010 -34 2012 -32
rect 1997 -35 2012 -34
rect 2017 -32 2021 -30
rect 2017 -34 2018 -32
rect 2020 -34 2021 -32
rect 2017 -39 2021 -34
rect 2040 -27 2044 -25
rect 2048 -21 2052 -10
rect 2048 -23 2054 -21
rect 2048 -25 2051 -23
rect 2053 -25 2054 -23
rect 2048 -27 2054 -25
rect 2048 -30 2052 -27
rect 2032 -34 2052 -30
rect 2032 -38 2036 -34
rect 1996 -40 2018 -39
rect 99 -45 100 -43
rect 102 -45 103 -43
rect 247 -45 248 -43
rect 250 -45 251 -43
rect 99 -48 103 -45
rect 155 -46 161 -45
rect 155 -48 157 -46
rect 159 -48 161 -46
rect 189 -46 195 -45
rect 189 -48 191 -46
rect 193 -48 195 -46
rect 247 -48 251 -45
rect 267 -45 273 -44
rect 267 -47 269 -45
rect 271 -47 273 -45
rect 267 -48 273 -47
rect 286 -45 292 -44
rect 286 -47 288 -45
rect 290 -47 292 -45
rect 286 -48 292 -47
rect 366 -45 367 -43
rect 369 -45 370 -43
rect 514 -45 515 -43
rect 517 -45 518 -43
rect 366 -48 370 -45
rect 422 -46 428 -45
rect 422 -48 424 -46
rect 426 -48 428 -46
rect 456 -46 462 -45
rect 456 -48 458 -46
rect 460 -48 462 -46
rect 514 -48 518 -45
rect 534 -45 540 -44
rect 534 -47 536 -45
rect 538 -47 540 -45
rect 534 -48 540 -47
rect 553 -45 559 -44
rect 553 -47 555 -45
rect 557 -47 559 -45
rect 553 -48 559 -47
rect 633 -45 634 -43
rect 636 -45 637 -43
rect 781 -45 782 -43
rect 784 -45 785 -43
rect 633 -48 637 -45
rect 689 -46 695 -45
rect 689 -48 691 -46
rect 693 -48 695 -46
rect 723 -46 729 -45
rect 723 -48 725 -46
rect 727 -48 729 -46
rect 781 -48 785 -45
rect 801 -45 807 -44
rect 801 -47 803 -45
rect 805 -47 807 -45
rect 801 -48 807 -47
rect 820 -45 826 -44
rect 820 -47 822 -45
rect 824 -47 826 -45
rect 820 -48 826 -47
rect 900 -45 901 -43
rect 903 -45 904 -43
rect 1048 -45 1049 -43
rect 1051 -45 1052 -43
rect 900 -48 904 -45
rect 956 -46 962 -45
rect 956 -48 958 -46
rect 960 -48 962 -46
rect 990 -46 996 -45
rect 990 -48 992 -46
rect 994 -48 996 -46
rect 1048 -48 1052 -45
rect 1068 -45 1074 -44
rect 1068 -47 1070 -45
rect 1072 -47 1074 -45
rect 1068 -48 1074 -47
rect 1087 -45 1093 -44
rect 1087 -47 1089 -45
rect 1091 -47 1093 -45
rect 1087 -48 1093 -47
rect 1167 -45 1168 -43
rect 1170 -45 1171 -43
rect 1315 -45 1316 -43
rect 1318 -45 1319 -43
rect 1167 -48 1171 -45
rect 1223 -46 1229 -45
rect 1223 -48 1225 -46
rect 1227 -48 1229 -46
rect 1257 -46 1263 -45
rect 1257 -48 1259 -46
rect 1261 -48 1263 -46
rect 1315 -48 1319 -45
rect 1335 -45 1341 -44
rect 1335 -47 1337 -45
rect 1339 -47 1341 -45
rect 1335 -48 1341 -47
rect 1354 -45 1360 -44
rect 1354 -47 1356 -45
rect 1358 -47 1360 -45
rect 1354 -48 1360 -47
rect 1434 -45 1435 -43
rect 1437 -45 1438 -43
rect 1582 -45 1583 -43
rect 1585 -45 1586 -43
rect 1434 -48 1438 -45
rect 1490 -46 1496 -45
rect 1490 -48 1492 -46
rect 1494 -48 1496 -46
rect 1524 -46 1530 -45
rect 1524 -48 1526 -46
rect 1528 -48 1530 -46
rect 1582 -48 1586 -45
rect 1602 -45 1608 -44
rect 1602 -47 1604 -45
rect 1606 -47 1608 -45
rect 1602 -48 1608 -47
rect 1621 -45 1627 -44
rect 1621 -47 1623 -45
rect 1625 -47 1627 -45
rect 1621 -48 1627 -47
rect 1701 -45 1702 -43
rect 1704 -45 1705 -43
rect 1849 -45 1850 -43
rect 1852 -45 1853 -43
rect 1701 -48 1705 -45
rect 1757 -46 1763 -45
rect 1757 -48 1759 -46
rect 1761 -48 1763 -46
rect 1791 -46 1797 -45
rect 1791 -48 1793 -46
rect 1795 -48 1797 -46
rect 1849 -48 1853 -45
rect 1869 -45 1875 -44
rect 1869 -47 1871 -45
rect 1873 -47 1875 -45
rect 1869 -48 1875 -47
rect 1888 -45 1894 -44
rect 1888 -47 1890 -45
rect 1892 -47 1894 -45
rect 1888 -48 1894 -47
rect 1926 -48 1932 -42
rect 1987 -43 1991 -41
rect 1996 -42 1998 -40
rect 2000 -41 2018 -40
rect 2020 -41 2021 -39
rect 2000 -42 2021 -41
rect 2026 -39 2036 -38
rect 2026 -41 2028 -39
rect 2030 -41 2036 -39
rect 2026 -42 2036 -41
rect 2087 -6 2091 -2
rect 2110 -6 2134 -2
rect 2074 -7 2114 -6
rect 2074 -9 2088 -7
rect 2090 -9 2114 -7
rect 2074 -10 2114 -9
rect 2074 -21 2078 -10
rect 2122 -11 2126 -9
rect 2130 -10 2136 -6
rect 2122 -13 2123 -11
rect 2125 -13 2126 -11
rect 2122 -14 2126 -13
rect 2122 -18 2129 -14
rect 2072 -23 2078 -21
rect 2072 -25 2073 -23
rect 2075 -25 2078 -23
rect 2072 -27 2078 -25
rect 2082 -23 2086 -18
rect 2082 -25 2083 -23
rect 2085 -25 2086 -23
rect 2082 -27 2086 -25
rect 2074 -30 2078 -27
rect 2074 -34 2094 -30
rect 2090 -38 2094 -34
rect 2125 -29 2129 -18
rect 2132 -20 2136 -10
rect 2132 -22 2133 -20
rect 2135 -22 2136 -20
rect 2132 -24 2136 -22
rect 2125 -30 2143 -29
rect 2105 -32 2109 -30
rect 2125 -31 2139 -30
rect 2105 -34 2106 -32
rect 2108 -34 2109 -32
rect 2090 -39 2100 -38
rect 2090 -41 2096 -39
rect 2098 -41 2100 -39
rect 2090 -42 2100 -41
rect 2105 -39 2109 -34
rect 2114 -32 2139 -31
rect 2141 -32 2143 -30
rect 2114 -34 2116 -32
rect 2118 -33 2143 -32
rect 2168 -6 2172 -2
rect 2168 -10 2183 -6
rect 2158 -19 2164 -18
rect 2118 -34 2129 -33
rect 2114 -35 2129 -34
rect 2179 -23 2183 -10
rect 2186 -13 2187 -2
rect 2226 -2 2239 -1
rect 2226 -4 2228 -2
rect 2230 -4 2239 -2
rect 2226 -5 2239 -4
rect 2235 -9 2251 -5
rect 2179 -25 2180 -23
rect 2182 -25 2183 -23
rect 2179 -31 2183 -25
rect 2223 -13 2227 -11
rect 2165 -32 2183 -31
rect 2165 -34 2167 -32
rect 2169 -34 2183 -32
rect 2165 -35 2183 -34
rect 2199 -14 2224 -13
rect 2199 -16 2201 -14
rect 2203 -15 2224 -14
rect 2226 -15 2227 -13
rect 2203 -16 2227 -15
rect 2199 -17 2227 -16
rect 2105 -41 2106 -39
rect 2108 -40 2130 -39
rect 2108 -41 2126 -40
rect 2105 -42 2126 -41
rect 2128 -42 2130 -40
rect 2199 -37 2203 -17
rect 2223 -27 2227 -17
rect 2243 -22 2244 -16
rect 2247 -26 2251 -9
rect 2223 -29 2234 -27
rect 2223 -31 2231 -29
rect 2233 -31 2234 -29
rect 2247 -28 2252 -26
rect 2247 -30 2249 -28
rect 2251 -30 2252 -28
rect 2223 -33 2234 -31
rect 2237 -32 2252 -30
rect 2237 -34 2251 -32
rect 2199 -38 2205 -37
rect 2199 -40 2201 -38
rect 2203 -40 2205 -38
rect 2199 -41 2205 -40
rect 2209 -38 2215 -37
rect 2209 -40 2211 -38
rect 2213 -40 2215 -38
rect 2237 -39 2241 -34
rect 2294 -2 2307 -1
rect 2294 -4 2296 -2
rect 2298 -4 2307 -2
rect 2294 -5 2307 -4
rect 2303 -9 2319 -5
rect 2291 -13 2295 -11
rect 1996 -43 2021 -42
rect 2105 -43 2130 -42
rect 2135 -43 2139 -41
rect 1987 -45 1988 -43
rect 1990 -45 1991 -43
rect 2135 -45 2136 -43
rect 2138 -45 2139 -43
rect 1987 -48 1991 -45
rect 2043 -46 2049 -45
rect 2043 -48 2045 -46
rect 2047 -48 2049 -46
rect 2077 -46 2083 -45
rect 2077 -48 2079 -46
rect 2081 -48 2083 -46
rect 2135 -48 2139 -45
rect 2155 -45 2161 -44
rect 2155 -47 2157 -45
rect 2159 -47 2161 -45
rect 2155 -48 2161 -47
rect 2174 -45 2180 -44
rect 2174 -47 2176 -45
rect 2178 -47 2180 -45
rect 2174 -48 2180 -47
rect 2209 -48 2215 -40
rect 2226 -40 2241 -39
rect 2226 -42 2228 -40
rect 2230 -42 2241 -40
rect 2226 -43 2241 -42
rect 2244 -40 2248 -38
rect 2244 -42 2245 -40
rect 2247 -42 2248 -40
rect 2267 -14 2292 -13
rect 2267 -16 2269 -14
rect 2271 -15 2292 -14
rect 2294 -15 2295 -13
rect 2271 -16 2295 -15
rect 2267 -17 2295 -16
rect 2267 -37 2271 -17
rect 2291 -27 2295 -17
rect 2311 -22 2312 -16
rect 2315 -26 2319 -9
rect 2291 -29 2302 -27
rect 2291 -31 2299 -29
rect 2301 -31 2302 -29
rect 2315 -28 2320 -26
rect 2315 -30 2317 -28
rect 2319 -30 2320 -28
rect 2291 -33 2302 -31
rect 2305 -32 2320 -30
rect 2305 -34 2319 -32
rect 2267 -38 2273 -37
rect 2267 -40 2269 -38
rect 2271 -40 2273 -38
rect 2267 -41 2273 -40
rect 2277 -38 2283 -37
rect 2277 -40 2279 -38
rect 2281 -40 2283 -38
rect 2305 -39 2309 -34
rect 2244 -48 2248 -42
rect 2277 -48 2283 -40
rect 2294 -40 2309 -39
rect 2294 -42 2296 -40
rect 2298 -42 2309 -40
rect 2294 -43 2309 -42
rect 2312 -40 2316 -38
rect 2312 -42 2313 -40
rect 2315 -42 2316 -40
rect 2312 -48 2316 -42
rect 99 -67 103 -64
rect 155 -66 157 -64
rect 159 -66 161 -64
rect 155 -67 161 -66
rect 189 -66 191 -64
rect 193 -66 195 -64
rect 189 -67 195 -66
rect 247 -67 251 -64
rect 99 -69 100 -67
rect 102 -69 103 -67
rect 247 -69 248 -67
rect 250 -69 251 -67
rect 267 -65 273 -64
rect 267 -67 269 -65
rect 271 -67 273 -65
rect 267 -68 273 -67
rect 286 -65 292 -64
rect 286 -67 288 -65
rect 290 -67 292 -65
rect 286 -68 292 -67
rect 366 -67 370 -64
rect 422 -66 424 -64
rect 426 -66 428 -64
rect 422 -67 428 -66
rect 456 -66 458 -64
rect 460 -66 462 -64
rect 456 -67 462 -66
rect 514 -67 518 -64
rect 366 -69 367 -67
rect 369 -69 370 -67
rect 514 -69 515 -67
rect 517 -69 518 -67
rect 534 -65 540 -64
rect 534 -67 536 -65
rect 538 -67 540 -65
rect 534 -68 540 -67
rect 553 -65 559 -64
rect 553 -67 555 -65
rect 557 -67 559 -65
rect 553 -68 559 -67
rect 633 -67 637 -64
rect 689 -66 691 -64
rect 693 -66 695 -64
rect 689 -67 695 -66
rect 723 -66 725 -64
rect 727 -66 729 -64
rect 723 -67 729 -66
rect 781 -67 785 -64
rect 633 -69 634 -67
rect 636 -69 637 -67
rect 781 -69 782 -67
rect 784 -69 785 -67
rect 801 -65 807 -64
rect 801 -67 803 -65
rect 805 -67 807 -65
rect 801 -68 807 -67
rect 820 -65 826 -64
rect 820 -67 822 -65
rect 824 -67 826 -65
rect 820 -68 826 -67
rect 900 -67 904 -64
rect 956 -66 958 -64
rect 960 -66 962 -64
rect 956 -67 962 -66
rect 990 -66 992 -64
rect 994 -66 996 -64
rect 990 -67 996 -66
rect 1048 -67 1052 -64
rect 900 -69 901 -67
rect 903 -69 904 -67
rect 1048 -69 1049 -67
rect 1051 -69 1052 -67
rect 1068 -65 1074 -64
rect 1068 -67 1070 -65
rect 1072 -67 1074 -65
rect 1068 -68 1074 -67
rect 1087 -65 1093 -64
rect 1087 -67 1089 -65
rect 1091 -67 1093 -65
rect 1087 -68 1093 -67
rect 1167 -67 1171 -64
rect 1223 -66 1225 -64
rect 1227 -66 1229 -64
rect 1223 -67 1229 -66
rect 1257 -66 1259 -64
rect 1261 -66 1263 -64
rect 1257 -67 1263 -66
rect 1315 -67 1319 -64
rect 1167 -69 1168 -67
rect 1170 -69 1171 -67
rect 1315 -69 1316 -67
rect 1318 -69 1319 -67
rect 1335 -65 1341 -64
rect 1335 -67 1337 -65
rect 1339 -67 1341 -65
rect 1335 -68 1341 -67
rect 1354 -65 1360 -64
rect 1354 -67 1356 -65
rect 1358 -67 1360 -65
rect 1354 -68 1360 -67
rect 1434 -67 1438 -64
rect 1490 -66 1492 -64
rect 1494 -66 1496 -64
rect 1490 -67 1496 -66
rect 1524 -66 1526 -64
rect 1528 -66 1530 -64
rect 1524 -67 1530 -66
rect 1582 -67 1586 -64
rect 1434 -69 1435 -67
rect 1437 -69 1438 -67
rect 1582 -69 1583 -67
rect 1585 -69 1586 -67
rect 1602 -65 1608 -64
rect 1602 -67 1604 -65
rect 1606 -67 1608 -65
rect 1602 -68 1608 -67
rect 1621 -65 1627 -64
rect 1621 -67 1623 -65
rect 1625 -67 1627 -65
rect 1621 -68 1627 -67
rect 1701 -67 1705 -64
rect 1757 -66 1759 -64
rect 1761 -66 1763 -64
rect 1757 -67 1763 -66
rect 1791 -66 1793 -64
rect 1795 -66 1797 -64
rect 1791 -67 1797 -66
rect 1849 -67 1853 -64
rect 1701 -69 1702 -67
rect 1704 -69 1705 -67
rect 1849 -69 1850 -67
rect 1852 -69 1853 -67
rect 1869 -65 1875 -64
rect 1869 -67 1871 -65
rect 1873 -67 1875 -65
rect 1869 -68 1875 -67
rect 1888 -65 1894 -64
rect 1888 -67 1890 -65
rect 1892 -67 1894 -65
rect 1888 -68 1894 -67
rect 8 -71 28 -70
rect 8 -73 10 -71
rect 12 -73 28 -71
rect 8 -74 28 -73
rect 24 -78 28 -74
rect 48 -71 68 -70
rect 48 -73 50 -71
rect 52 -73 68 -71
rect 48 -74 68 -73
rect 39 -77 40 -75
rect 24 -82 36 -78
rect 32 -87 36 -82
rect 32 -89 33 -87
rect 35 -89 36 -87
rect 32 -101 36 -89
rect 64 -78 68 -74
rect 79 -77 80 -75
rect 64 -82 76 -78
rect 72 -87 76 -82
rect 72 -89 73 -87
rect 75 -89 76 -87
rect 19 -104 36 -101
rect 19 -106 20 -104
rect 22 -105 36 -104
rect 22 -106 23 -105
rect 8 -111 14 -110
rect 8 -113 10 -111
rect 12 -113 14 -111
rect 8 -120 14 -113
rect 19 -111 23 -106
rect 72 -101 76 -89
rect 59 -104 76 -101
rect 59 -106 60 -104
rect 62 -105 76 -104
rect 62 -106 63 -105
rect 19 -113 20 -111
rect 22 -113 23 -111
rect 19 -115 23 -113
rect 28 -109 34 -108
rect 28 -111 30 -109
rect 32 -111 34 -109
rect 28 -120 34 -111
rect 48 -111 54 -110
rect 48 -113 50 -111
rect 52 -113 54 -111
rect 48 -120 54 -113
rect 59 -111 63 -106
rect 99 -71 103 -69
rect 108 -70 133 -69
rect 217 -70 242 -69
rect 108 -72 110 -70
rect 112 -71 133 -70
rect 112 -72 130 -71
rect 108 -73 130 -72
rect 132 -73 133 -71
rect 109 -78 124 -77
rect 109 -79 120 -78
rect 95 -80 120 -79
rect 122 -80 124 -78
rect 95 -82 97 -80
rect 99 -81 124 -80
rect 129 -78 133 -73
rect 138 -71 148 -70
rect 138 -73 140 -71
rect 142 -73 148 -71
rect 138 -74 148 -73
rect 129 -80 130 -78
rect 132 -80 133 -78
rect 99 -82 113 -81
rect 129 -82 133 -80
rect 95 -83 113 -82
rect 102 -90 106 -88
rect 102 -92 103 -90
rect 105 -92 106 -90
rect 102 -102 106 -92
rect 109 -94 113 -83
rect 144 -78 148 -74
rect 144 -82 164 -78
rect 160 -85 164 -82
rect 152 -87 156 -85
rect 152 -89 153 -87
rect 155 -89 156 -87
rect 152 -94 156 -89
rect 160 -87 166 -85
rect 160 -89 163 -87
rect 165 -89 166 -87
rect 160 -91 166 -89
rect 109 -98 116 -94
rect 112 -99 116 -98
rect 112 -101 113 -99
rect 115 -101 116 -99
rect 102 -106 108 -102
rect 112 -103 116 -101
rect 160 -102 164 -91
rect 124 -103 164 -102
rect 124 -105 148 -103
rect 150 -105 164 -103
rect 124 -106 164 -105
rect 59 -113 60 -111
rect 62 -113 63 -111
rect 59 -115 63 -113
rect 68 -109 74 -108
rect 68 -111 70 -109
rect 72 -111 74 -109
rect 104 -110 128 -106
rect 147 -110 151 -106
rect 202 -71 212 -70
rect 202 -73 208 -71
rect 210 -73 212 -71
rect 202 -74 212 -73
rect 217 -71 238 -70
rect 217 -73 218 -71
rect 220 -72 238 -71
rect 240 -72 242 -70
rect 247 -71 251 -69
rect 220 -73 242 -72
rect 202 -78 206 -74
rect 186 -82 206 -78
rect 186 -85 190 -82
rect 184 -87 190 -85
rect 184 -89 185 -87
rect 187 -89 190 -87
rect 184 -91 190 -89
rect 186 -102 190 -91
rect 194 -87 198 -85
rect 217 -78 221 -73
rect 315 -71 335 -70
rect 315 -73 317 -71
rect 319 -73 335 -71
rect 315 -74 335 -73
rect 217 -80 218 -78
rect 220 -80 221 -78
rect 217 -82 221 -80
rect 226 -78 241 -77
rect 226 -80 228 -78
rect 230 -79 241 -78
rect 230 -80 255 -79
rect 226 -81 251 -80
rect 237 -82 251 -81
rect 253 -82 255 -80
rect 237 -83 255 -82
rect 194 -89 195 -87
rect 197 -89 198 -87
rect 194 -94 198 -89
rect 237 -94 241 -83
rect 234 -98 241 -94
rect 244 -90 248 -88
rect 244 -92 245 -90
rect 247 -92 248 -90
rect 234 -99 238 -98
rect 234 -101 235 -99
rect 237 -101 238 -99
rect 186 -103 226 -102
rect 234 -103 238 -101
rect 244 -102 248 -92
rect 277 -78 295 -77
rect 277 -80 279 -78
rect 281 -80 295 -78
rect 277 -81 295 -80
rect 291 -87 295 -81
rect 291 -89 292 -87
rect 294 -89 295 -87
rect 270 -94 276 -93
rect 186 -105 200 -103
rect 202 -105 226 -103
rect 186 -106 226 -105
rect 242 -106 248 -102
rect 199 -110 203 -106
rect 222 -110 246 -106
rect 291 -102 295 -89
rect 280 -106 295 -102
rect 280 -110 284 -106
rect 298 -110 299 -99
rect 331 -78 335 -74
rect 346 -77 347 -75
rect 331 -82 343 -78
rect 339 -87 343 -82
rect 339 -89 340 -87
rect 342 -89 343 -87
rect 339 -101 343 -89
rect 326 -104 343 -101
rect 326 -106 327 -104
rect 329 -105 343 -104
rect 329 -106 330 -105
rect 68 -120 74 -111
rect 134 -111 140 -110
rect 134 -113 136 -111
rect 138 -113 140 -111
rect 99 -118 105 -117
rect 99 -120 101 -118
rect 103 -120 105 -118
rect 134 -118 140 -113
rect 147 -112 148 -110
rect 150 -112 151 -110
rect 147 -114 151 -112
rect 156 -111 162 -110
rect 156 -113 158 -111
rect 160 -113 162 -111
rect 134 -120 136 -118
rect 138 -120 140 -118
rect 156 -118 162 -113
rect 156 -120 158 -118
rect 160 -120 162 -118
rect 188 -111 194 -110
rect 188 -113 190 -111
rect 192 -113 194 -111
rect 188 -118 194 -113
rect 199 -112 200 -110
rect 202 -112 203 -110
rect 199 -114 203 -112
rect 210 -111 216 -110
rect 210 -113 212 -111
rect 214 -113 216 -111
rect 188 -120 190 -118
rect 192 -120 194 -118
rect 210 -118 216 -113
rect 267 -111 284 -110
rect 267 -113 269 -111
rect 271 -113 284 -111
rect 267 -114 284 -113
rect 315 -111 321 -110
rect 315 -113 317 -111
rect 319 -113 321 -111
rect 210 -120 212 -118
rect 214 -120 216 -118
rect 245 -118 251 -117
rect 245 -120 247 -118
rect 249 -120 251 -118
rect 286 -118 292 -117
rect 286 -120 288 -118
rect 290 -120 292 -118
rect 315 -120 321 -113
rect 326 -111 330 -106
rect 366 -71 370 -69
rect 375 -70 400 -69
rect 484 -70 509 -69
rect 375 -72 377 -70
rect 379 -71 400 -70
rect 379 -72 397 -71
rect 375 -73 397 -72
rect 399 -73 400 -71
rect 376 -78 391 -77
rect 376 -79 387 -78
rect 362 -80 387 -79
rect 389 -80 391 -78
rect 362 -82 364 -80
rect 366 -81 391 -80
rect 396 -78 400 -73
rect 405 -71 415 -70
rect 405 -73 407 -71
rect 409 -73 415 -71
rect 405 -74 415 -73
rect 396 -80 397 -78
rect 399 -80 400 -78
rect 366 -82 380 -81
rect 396 -82 400 -80
rect 362 -83 380 -82
rect 369 -90 373 -88
rect 369 -92 370 -90
rect 372 -92 373 -90
rect 369 -102 373 -92
rect 376 -94 380 -83
rect 411 -78 415 -74
rect 411 -82 431 -78
rect 427 -85 431 -82
rect 419 -87 423 -85
rect 419 -89 420 -87
rect 422 -89 423 -87
rect 419 -94 423 -89
rect 427 -87 433 -85
rect 427 -89 430 -87
rect 432 -89 433 -87
rect 427 -91 433 -89
rect 376 -98 383 -94
rect 379 -99 383 -98
rect 379 -101 380 -99
rect 382 -101 383 -99
rect 369 -106 375 -102
rect 379 -103 383 -101
rect 427 -102 431 -91
rect 391 -103 431 -102
rect 391 -105 415 -103
rect 417 -105 431 -103
rect 391 -106 431 -105
rect 326 -113 327 -111
rect 329 -113 330 -111
rect 326 -115 330 -113
rect 335 -109 341 -108
rect 335 -111 337 -109
rect 339 -111 341 -109
rect 371 -110 395 -106
rect 414 -110 418 -106
rect 469 -71 479 -70
rect 469 -73 475 -71
rect 477 -73 479 -71
rect 469 -74 479 -73
rect 484 -71 505 -70
rect 484 -73 485 -71
rect 487 -72 505 -71
rect 507 -72 509 -70
rect 514 -71 518 -69
rect 487 -73 509 -72
rect 469 -78 473 -74
rect 453 -82 473 -78
rect 453 -85 457 -82
rect 451 -87 457 -85
rect 451 -89 452 -87
rect 454 -89 457 -87
rect 451 -91 457 -89
rect 453 -102 457 -91
rect 461 -87 465 -85
rect 484 -78 488 -73
rect 582 -71 602 -70
rect 582 -73 584 -71
rect 586 -73 602 -71
rect 582 -74 602 -73
rect 484 -80 485 -78
rect 487 -80 488 -78
rect 484 -82 488 -80
rect 493 -78 508 -77
rect 493 -80 495 -78
rect 497 -79 508 -78
rect 497 -80 522 -79
rect 493 -81 518 -80
rect 504 -82 518 -81
rect 520 -82 522 -80
rect 504 -83 522 -82
rect 461 -89 462 -87
rect 464 -89 465 -87
rect 461 -94 465 -89
rect 504 -94 508 -83
rect 501 -98 508 -94
rect 511 -90 515 -88
rect 511 -92 512 -90
rect 514 -92 515 -90
rect 501 -99 505 -98
rect 501 -101 502 -99
rect 504 -101 505 -99
rect 453 -103 493 -102
rect 501 -103 505 -101
rect 511 -102 515 -92
rect 544 -78 562 -77
rect 544 -80 546 -78
rect 548 -80 562 -78
rect 544 -81 562 -80
rect 558 -87 562 -81
rect 558 -89 559 -87
rect 561 -89 562 -87
rect 537 -94 543 -93
rect 453 -105 467 -103
rect 469 -105 493 -103
rect 453 -106 493 -105
rect 509 -106 515 -102
rect 466 -110 470 -106
rect 489 -110 513 -106
rect 558 -102 562 -89
rect 547 -106 562 -102
rect 547 -110 551 -106
rect 565 -110 566 -99
rect 598 -78 602 -74
rect 613 -77 614 -75
rect 598 -82 610 -78
rect 606 -87 610 -82
rect 606 -89 607 -87
rect 609 -89 610 -87
rect 606 -101 610 -89
rect 593 -104 610 -101
rect 593 -106 594 -104
rect 596 -105 610 -104
rect 596 -106 597 -105
rect 335 -120 341 -111
rect 401 -111 407 -110
rect 401 -113 403 -111
rect 405 -113 407 -111
rect 366 -118 372 -117
rect 366 -120 368 -118
rect 370 -120 372 -118
rect 401 -118 407 -113
rect 414 -112 415 -110
rect 417 -112 418 -110
rect 414 -114 418 -112
rect 423 -111 429 -110
rect 423 -113 425 -111
rect 427 -113 429 -111
rect 401 -120 403 -118
rect 405 -120 407 -118
rect 423 -118 429 -113
rect 423 -120 425 -118
rect 427 -120 429 -118
rect 455 -111 461 -110
rect 455 -113 457 -111
rect 459 -113 461 -111
rect 455 -118 461 -113
rect 466 -112 467 -110
rect 469 -112 470 -110
rect 466 -114 470 -112
rect 477 -111 483 -110
rect 477 -113 479 -111
rect 481 -113 483 -111
rect 455 -120 457 -118
rect 459 -120 461 -118
rect 477 -118 483 -113
rect 534 -111 551 -110
rect 534 -113 536 -111
rect 538 -113 551 -111
rect 534 -114 551 -113
rect 582 -111 588 -110
rect 582 -113 584 -111
rect 586 -113 588 -111
rect 477 -120 479 -118
rect 481 -120 483 -118
rect 512 -118 518 -117
rect 512 -120 514 -118
rect 516 -120 518 -118
rect 553 -118 559 -117
rect 553 -120 555 -118
rect 557 -120 559 -118
rect 582 -120 588 -113
rect 593 -111 597 -106
rect 633 -71 637 -69
rect 642 -70 667 -69
rect 751 -70 776 -69
rect 642 -72 644 -70
rect 646 -71 667 -70
rect 646 -72 664 -71
rect 642 -73 664 -72
rect 666 -73 667 -71
rect 643 -78 658 -77
rect 643 -79 654 -78
rect 629 -80 654 -79
rect 656 -80 658 -78
rect 629 -82 631 -80
rect 633 -81 658 -80
rect 663 -78 667 -73
rect 672 -71 682 -70
rect 672 -73 674 -71
rect 676 -73 682 -71
rect 672 -74 682 -73
rect 663 -80 664 -78
rect 666 -80 667 -78
rect 633 -82 647 -81
rect 663 -82 667 -80
rect 629 -83 647 -82
rect 636 -90 640 -88
rect 636 -92 637 -90
rect 639 -92 640 -90
rect 636 -102 640 -92
rect 643 -94 647 -83
rect 678 -78 682 -74
rect 678 -82 698 -78
rect 694 -85 698 -82
rect 686 -87 690 -85
rect 686 -89 687 -87
rect 689 -89 690 -87
rect 686 -94 690 -89
rect 694 -87 700 -85
rect 694 -89 697 -87
rect 699 -89 700 -87
rect 694 -91 700 -89
rect 643 -98 650 -94
rect 646 -99 650 -98
rect 646 -101 647 -99
rect 649 -101 650 -99
rect 636 -106 642 -102
rect 646 -103 650 -101
rect 694 -102 698 -91
rect 658 -103 698 -102
rect 658 -105 682 -103
rect 684 -105 698 -103
rect 658 -106 698 -105
rect 593 -113 594 -111
rect 596 -113 597 -111
rect 593 -115 597 -113
rect 602 -109 608 -108
rect 602 -111 604 -109
rect 606 -111 608 -109
rect 638 -110 662 -106
rect 681 -110 685 -106
rect 736 -71 746 -70
rect 736 -73 742 -71
rect 744 -73 746 -71
rect 736 -74 746 -73
rect 751 -71 772 -70
rect 751 -73 752 -71
rect 754 -72 772 -71
rect 774 -72 776 -70
rect 781 -71 785 -69
rect 754 -73 776 -72
rect 736 -78 740 -74
rect 720 -82 740 -78
rect 720 -85 724 -82
rect 718 -87 724 -85
rect 718 -89 719 -87
rect 721 -89 724 -87
rect 718 -91 724 -89
rect 720 -102 724 -91
rect 728 -87 732 -85
rect 751 -78 755 -73
rect 849 -71 869 -70
rect 849 -73 851 -71
rect 853 -73 869 -71
rect 849 -74 869 -73
rect 751 -80 752 -78
rect 754 -80 755 -78
rect 751 -82 755 -80
rect 760 -78 775 -77
rect 760 -80 762 -78
rect 764 -79 775 -78
rect 764 -80 789 -79
rect 760 -81 785 -80
rect 771 -82 785 -81
rect 787 -82 789 -80
rect 771 -83 789 -82
rect 728 -89 729 -87
rect 731 -89 732 -87
rect 728 -94 732 -89
rect 771 -94 775 -83
rect 768 -98 775 -94
rect 778 -90 782 -88
rect 778 -92 779 -90
rect 781 -92 782 -90
rect 768 -99 772 -98
rect 768 -101 769 -99
rect 771 -101 772 -99
rect 720 -103 760 -102
rect 768 -103 772 -101
rect 778 -102 782 -92
rect 811 -78 829 -77
rect 811 -80 813 -78
rect 815 -80 829 -78
rect 811 -81 829 -80
rect 825 -87 829 -81
rect 825 -89 826 -87
rect 828 -89 829 -87
rect 804 -94 810 -93
rect 720 -105 734 -103
rect 736 -105 760 -103
rect 720 -106 760 -105
rect 776 -106 782 -102
rect 733 -110 737 -106
rect 756 -110 780 -106
rect 825 -102 829 -89
rect 814 -106 829 -102
rect 814 -110 818 -106
rect 832 -110 833 -99
rect 865 -78 869 -74
rect 880 -77 881 -75
rect 865 -82 877 -78
rect 873 -87 877 -82
rect 873 -89 874 -87
rect 876 -89 877 -87
rect 873 -101 877 -89
rect 860 -104 877 -101
rect 860 -106 861 -104
rect 863 -105 877 -104
rect 863 -106 864 -105
rect 602 -120 608 -111
rect 668 -111 674 -110
rect 668 -113 670 -111
rect 672 -113 674 -111
rect 633 -118 639 -117
rect 633 -120 635 -118
rect 637 -120 639 -118
rect 668 -118 674 -113
rect 681 -112 682 -110
rect 684 -112 685 -110
rect 681 -114 685 -112
rect 690 -111 696 -110
rect 690 -113 692 -111
rect 694 -113 696 -111
rect 668 -120 670 -118
rect 672 -120 674 -118
rect 690 -118 696 -113
rect 690 -120 692 -118
rect 694 -120 696 -118
rect 722 -111 728 -110
rect 722 -113 724 -111
rect 726 -113 728 -111
rect 722 -118 728 -113
rect 733 -112 734 -110
rect 736 -112 737 -110
rect 733 -114 737 -112
rect 744 -111 750 -110
rect 744 -113 746 -111
rect 748 -113 750 -111
rect 722 -120 724 -118
rect 726 -120 728 -118
rect 744 -118 750 -113
rect 801 -111 818 -110
rect 801 -113 803 -111
rect 805 -113 818 -111
rect 801 -114 818 -113
rect 849 -111 855 -110
rect 849 -113 851 -111
rect 853 -113 855 -111
rect 744 -120 746 -118
rect 748 -120 750 -118
rect 779 -118 785 -117
rect 779 -120 781 -118
rect 783 -120 785 -118
rect 820 -118 826 -117
rect 820 -120 822 -118
rect 824 -120 826 -118
rect 849 -120 855 -113
rect 860 -111 864 -106
rect 900 -71 904 -69
rect 909 -70 934 -69
rect 1018 -70 1043 -69
rect 909 -72 911 -70
rect 913 -71 934 -70
rect 913 -72 931 -71
rect 909 -73 931 -72
rect 933 -73 934 -71
rect 910 -78 925 -77
rect 910 -79 921 -78
rect 896 -80 921 -79
rect 923 -80 925 -78
rect 896 -82 898 -80
rect 900 -81 925 -80
rect 930 -78 934 -73
rect 939 -71 949 -70
rect 939 -73 941 -71
rect 943 -73 949 -71
rect 939 -74 949 -73
rect 930 -80 931 -78
rect 933 -80 934 -78
rect 900 -82 914 -81
rect 930 -82 934 -80
rect 896 -83 914 -82
rect 903 -90 907 -88
rect 903 -92 904 -90
rect 906 -92 907 -90
rect 903 -102 907 -92
rect 910 -94 914 -83
rect 945 -78 949 -74
rect 945 -82 965 -78
rect 961 -85 965 -82
rect 953 -87 957 -85
rect 953 -89 954 -87
rect 956 -89 957 -87
rect 953 -94 957 -89
rect 961 -87 967 -85
rect 961 -89 964 -87
rect 966 -89 967 -87
rect 961 -91 967 -89
rect 910 -98 917 -94
rect 913 -99 917 -98
rect 913 -101 914 -99
rect 916 -101 917 -99
rect 903 -106 909 -102
rect 913 -103 917 -101
rect 961 -102 965 -91
rect 925 -103 965 -102
rect 925 -105 949 -103
rect 951 -105 965 -103
rect 925 -106 965 -105
rect 860 -113 861 -111
rect 863 -113 864 -111
rect 860 -115 864 -113
rect 869 -109 875 -108
rect 869 -111 871 -109
rect 873 -111 875 -109
rect 905 -110 929 -106
rect 948 -110 952 -106
rect 1003 -71 1013 -70
rect 1003 -73 1009 -71
rect 1011 -73 1013 -71
rect 1003 -74 1013 -73
rect 1018 -71 1039 -70
rect 1018 -73 1019 -71
rect 1021 -72 1039 -71
rect 1041 -72 1043 -70
rect 1048 -71 1052 -69
rect 1021 -73 1043 -72
rect 1003 -78 1007 -74
rect 987 -82 1007 -78
rect 987 -85 991 -82
rect 985 -87 991 -85
rect 985 -89 986 -87
rect 988 -89 991 -87
rect 985 -91 991 -89
rect 987 -102 991 -91
rect 995 -87 999 -85
rect 1018 -78 1022 -73
rect 1116 -71 1136 -70
rect 1116 -73 1118 -71
rect 1120 -73 1136 -71
rect 1116 -74 1136 -73
rect 1018 -80 1019 -78
rect 1021 -80 1022 -78
rect 1018 -82 1022 -80
rect 1027 -78 1042 -77
rect 1027 -80 1029 -78
rect 1031 -79 1042 -78
rect 1031 -80 1056 -79
rect 1027 -81 1052 -80
rect 1038 -82 1052 -81
rect 1054 -82 1056 -80
rect 1038 -83 1056 -82
rect 995 -89 996 -87
rect 998 -89 999 -87
rect 995 -94 999 -89
rect 1038 -94 1042 -83
rect 1035 -98 1042 -94
rect 1045 -90 1049 -88
rect 1045 -92 1046 -90
rect 1048 -92 1049 -90
rect 1035 -99 1039 -98
rect 1035 -101 1036 -99
rect 1038 -101 1039 -99
rect 987 -103 1027 -102
rect 1035 -103 1039 -101
rect 1045 -102 1049 -92
rect 1078 -78 1096 -77
rect 1078 -80 1080 -78
rect 1082 -80 1096 -78
rect 1078 -81 1096 -80
rect 1092 -87 1096 -81
rect 1092 -89 1093 -87
rect 1095 -89 1096 -87
rect 1071 -94 1077 -93
rect 987 -105 1001 -103
rect 1003 -105 1027 -103
rect 987 -106 1027 -105
rect 1043 -106 1049 -102
rect 1000 -110 1004 -106
rect 1023 -110 1047 -106
rect 1092 -102 1096 -89
rect 1081 -106 1096 -102
rect 1081 -110 1085 -106
rect 1099 -110 1100 -99
rect 1132 -78 1136 -74
rect 1147 -77 1148 -75
rect 1132 -82 1144 -78
rect 1140 -87 1144 -82
rect 1140 -89 1141 -87
rect 1143 -89 1144 -87
rect 1140 -101 1144 -89
rect 1127 -104 1144 -101
rect 1127 -106 1128 -104
rect 1130 -105 1144 -104
rect 1130 -106 1131 -105
rect 869 -120 875 -111
rect 935 -111 941 -110
rect 935 -113 937 -111
rect 939 -113 941 -111
rect 900 -118 906 -117
rect 900 -120 902 -118
rect 904 -120 906 -118
rect 935 -118 941 -113
rect 948 -112 949 -110
rect 951 -112 952 -110
rect 948 -114 952 -112
rect 957 -111 963 -110
rect 957 -113 959 -111
rect 961 -113 963 -111
rect 935 -120 937 -118
rect 939 -120 941 -118
rect 957 -118 963 -113
rect 957 -120 959 -118
rect 961 -120 963 -118
rect 989 -111 995 -110
rect 989 -113 991 -111
rect 993 -113 995 -111
rect 989 -118 995 -113
rect 1000 -112 1001 -110
rect 1003 -112 1004 -110
rect 1000 -114 1004 -112
rect 1011 -111 1017 -110
rect 1011 -113 1013 -111
rect 1015 -113 1017 -111
rect 989 -120 991 -118
rect 993 -120 995 -118
rect 1011 -118 1017 -113
rect 1068 -111 1085 -110
rect 1068 -113 1070 -111
rect 1072 -113 1085 -111
rect 1068 -114 1085 -113
rect 1116 -111 1122 -110
rect 1116 -113 1118 -111
rect 1120 -113 1122 -111
rect 1011 -120 1013 -118
rect 1015 -120 1017 -118
rect 1046 -118 1052 -117
rect 1046 -120 1048 -118
rect 1050 -120 1052 -118
rect 1087 -118 1093 -117
rect 1087 -120 1089 -118
rect 1091 -120 1093 -118
rect 1116 -120 1122 -113
rect 1127 -111 1131 -106
rect 1167 -71 1171 -69
rect 1176 -70 1201 -69
rect 1285 -70 1310 -69
rect 1176 -72 1178 -70
rect 1180 -71 1201 -70
rect 1180 -72 1198 -71
rect 1176 -73 1198 -72
rect 1200 -73 1201 -71
rect 1177 -78 1192 -77
rect 1177 -79 1188 -78
rect 1163 -80 1188 -79
rect 1190 -80 1192 -78
rect 1163 -82 1165 -80
rect 1167 -81 1192 -80
rect 1197 -78 1201 -73
rect 1206 -71 1216 -70
rect 1206 -73 1208 -71
rect 1210 -73 1216 -71
rect 1206 -74 1216 -73
rect 1197 -80 1198 -78
rect 1200 -80 1201 -78
rect 1167 -82 1181 -81
rect 1197 -82 1201 -80
rect 1163 -83 1181 -82
rect 1170 -90 1174 -88
rect 1170 -92 1171 -90
rect 1173 -92 1174 -90
rect 1170 -102 1174 -92
rect 1177 -94 1181 -83
rect 1212 -78 1216 -74
rect 1212 -82 1232 -78
rect 1228 -85 1232 -82
rect 1220 -87 1224 -85
rect 1220 -89 1221 -87
rect 1223 -89 1224 -87
rect 1220 -94 1224 -89
rect 1228 -87 1234 -85
rect 1228 -89 1231 -87
rect 1233 -89 1234 -87
rect 1228 -91 1234 -89
rect 1177 -98 1184 -94
rect 1180 -99 1184 -98
rect 1180 -101 1181 -99
rect 1183 -101 1184 -99
rect 1170 -106 1176 -102
rect 1180 -103 1184 -101
rect 1228 -102 1232 -91
rect 1192 -103 1232 -102
rect 1192 -105 1216 -103
rect 1218 -105 1232 -103
rect 1192 -106 1232 -105
rect 1127 -113 1128 -111
rect 1130 -113 1131 -111
rect 1127 -115 1131 -113
rect 1136 -109 1142 -108
rect 1136 -111 1138 -109
rect 1140 -111 1142 -109
rect 1172 -110 1196 -106
rect 1215 -110 1219 -106
rect 1270 -71 1280 -70
rect 1270 -73 1276 -71
rect 1278 -73 1280 -71
rect 1270 -74 1280 -73
rect 1285 -71 1306 -70
rect 1285 -73 1286 -71
rect 1288 -72 1306 -71
rect 1308 -72 1310 -70
rect 1315 -71 1319 -69
rect 1288 -73 1310 -72
rect 1270 -78 1274 -74
rect 1254 -82 1274 -78
rect 1254 -85 1258 -82
rect 1252 -87 1258 -85
rect 1252 -89 1253 -87
rect 1255 -89 1258 -87
rect 1252 -91 1258 -89
rect 1254 -102 1258 -91
rect 1262 -87 1266 -85
rect 1285 -78 1289 -73
rect 1383 -71 1403 -70
rect 1383 -73 1385 -71
rect 1387 -73 1403 -71
rect 1383 -74 1403 -73
rect 1285 -80 1286 -78
rect 1288 -80 1289 -78
rect 1285 -82 1289 -80
rect 1294 -78 1309 -77
rect 1294 -80 1296 -78
rect 1298 -79 1309 -78
rect 1298 -80 1323 -79
rect 1294 -81 1319 -80
rect 1305 -82 1319 -81
rect 1321 -82 1323 -80
rect 1305 -83 1323 -82
rect 1262 -89 1263 -87
rect 1265 -89 1266 -87
rect 1262 -94 1266 -89
rect 1305 -94 1309 -83
rect 1302 -98 1309 -94
rect 1312 -90 1316 -88
rect 1312 -92 1313 -90
rect 1315 -92 1316 -90
rect 1302 -99 1306 -98
rect 1302 -101 1303 -99
rect 1305 -101 1306 -99
rect 1254 -103 1294 -102
rect 1302 -103 1306 -101
rect 1312 -102 1316 -92
rect 1345 -78 1363 -77
rect 1345 -80 1347 -78
rect 1349 -80 1363 -78
rect 1345 -81 1363 -80
rect 1359 -87 1363 -81
rect 1359 -89 1360 -87
rect 1362 -89 1363 -87
rect 1338 -94 1344 -93
rect 1254 -105 1268 -103
rect 1270 -105 1294 -103
rect 1254 -106 1294 -105
rect 1310 -106 1316 -102
rect 1267 -110 1271 -106
rect 1290 -110 1314 -106
rect 1359 -102 1363 -89
rect 1348 -106 1363 -102
rect 1348 -110 1352 -106
rect 1366 -110 1367 -99
rect 1399 -78 1403 -74
rect 1414 -77 1415 -75
rect 1399 -82 1411 -78
rect 1407 -87 1411 -82
rect 1407 -89 1408 -87
rect 1410 -89 1411 -87
rect 1407 -101 1411 -89
rect 1394 -104 1411 -101
rect 1394 -106 1395 -104
rect 1397 -105 1411 -104
rect 1397 -106 1398 -105
rect 1136 -120 1142 -111
rect 1202 -111 1208 -110
rect 1202 -113 1204 -111
rect 1206 -113 1208 -111
rect 1167 -118 1173 -117
rect 1167 -120 1169 -118
rect 1171 -120 1173 -118
rect 1202 -118 1208 -113
rect 1215 -112 1216 -110
rect 1218 -112 1219 -110
rect 1215 -114 1219 -112
rect 1224 -111 1230 -110
rect 1224 -113 1226 -111
rect 1228 -113 1230 -111
rect 1202 -120 1204 -118
rect 1206 -120 1208 -118
rect 1224 -118 1230 -113
rect 1224 -120 1226 -118
rect 1228 -120 1230 -118
rect 1256 -111 1262 -110
rect 1256 -113 1258 -111
rect 1260 -113 1262 -111
rect 1256 -118 1262 -113
rect 1267 -112 1268 -110
rect 1270 -112 1271 -110
rect 1267 -114 1271 -112
rect 1278 -111 1284 -110
rect 1278 -113 1280 -111
rect 1282 -113 1284 -111
rect 1256 -120 1258 -118
rect 1260 -120 1262 -118
rect 1278 -118 1284 -113
rect 1335 -111 1352 -110
rect 1335 -113 1337 -111
rect 1339 -113 1352 -111
rect 1335 -114 1352 -113
rect 1383 -111 1389 -110
rect 1383 -113 1385 -111
rect 1387 -113 1389 -111
rect 1278 -120 1280 -118
rect 1282 -120 1284 -118
rect 1313 -118 1319 -117
rect 1313 -120 1315 -118
rect 1317 -120 1319 -118
rect 1354 -118 1360 -117
rect 1354 -120 1356 -118
rect 1358 -120 1360 -118
rect 1383 -120 1389 -113
rect 1394 -111 1398 -106
rect 1434 -71 1438 -69
rect 1443 -70 1468 -69
rect 1552 -70 1577 -69
rect 1443 -72 1445 -70
rect 1447 -71 1468 -70
rect 1447 -72 1465 -71
rect 1443 -73 1465 -72
rect 1467 -73 1468 -71
rect 1444 -78 1459 -77
rect 1444 -79 1455 -78
rect 1430 -80 1455 -79
rect 1457 -80 1459 -78
rect 1430 -82 1432 -80
rect 1434 -81 1459 -80
rect 1464 -78 1468 -73
rect 1473 -71 1483 -70
rect 1473 -73 1475 -71
rect 1477 -73 1483 -71
rect 1473 -74 1483 -73
rect 1464 -80 1465 -78
rect 1467 -80 1468 -78
rect 1434 -82 1448 -81
rect 1464 -82 1468 -80
rect 1430 -83 1448 -82
rect 1437 -90 1441 -88
rect 1437 -92 1438 -90
rect 1440 -92 1441 -90
rect 1437 -102 1441 -92
rect 1444 -94 1448 -83
rect 1479 -78 1483 -74
rect 1479 -82 1499 -78
rect 1495 -85 1499 -82
rect 1487 -87 1491 -85
rect 1487 -89 1488 -87
rect 1490 -89 1491 -87
rect 1487 -94 1491 -89
rect 1495 -87 1501 -85
rect 1495 -89 1498 -87
rect 1500 -89 1501 -87
rect 1495 -91 1501 -89
rect 1444 -98 1451 -94
rect 1447 -99 1451 -98
rect 1447 -101 1448 -99
rect 1450 -101 1451 -99
rect 1437 -106 1443 -102
rect 1447 -103 1451 -101
rect 1495 -102 1499 -91
rect 1459 -103 1499 -102
rect 1459 -105 1483 -103
rect 1485 -105 1499 -103
rect 1459 -106 1499 -105
rect 1394 -113 1395 -111
rect 1397 -113 1398 -111
rect 1394 -115 1398 -113
rect 1403 -109 1409 -108
rect 1403 -111 1405 -109
rect 1407 -111 1409 -109
rect 1439 -110 1463 -106
rect 1482 -110 1486 -106
rect 1537 -71 1547 -70
rect 1537 -73 1543 -71
rect 1545 -73 1547 -71
rect 1537 -74 1547 -73
rect 1552 -71 1573 -70
rect 1552 -73 1553 -71
rect 1555 -72 1573 -71
rect 1575 -72 1577 -70
rect 1582 -71 1586 -69
rect 1555 -73 1577 -72
rect 1537 -78 1541 -74
rect 1521 -82 1541 -78
rect 1521 -85 1525 -82
rect 1519 -87 1525 -85
rect 1519 -89 1520 -87
rect 1522 -89 1525 -87
rect 1519 -91 1525 -89
rect 1521 -102 1525 -91
rect 1529 -87 1533 -85
rect 1552 -78 1556 -73
rect 1650 -71 1670 -70
rect 1650 -73 1652 -71
rect 1654 -73 1670 -71
rect 1650 -74 1670 -73
rect 1552 -80 1553 -78
rect 1555 -80 1556 -78
rect 1552 -82 1556 -80
rect 1561 -78 1576 -77
rect 1561 -80 1563 -78
rect 1565 -79 1576 -78
rect 1565 -80 1590 -79
rect 1561 -81 1586 -80
rect 1572 -82 1586 -81
rect 1588 -82 1590 -80
rect 1572 -83 1590 -82
rect 1529 -89 1530 -87
rect 1532 -89 1533 -87
rect 1529 -94 1533 -89
rect 1572 -94 1576 -83
rect 1569 -98 1576 -94
rect 1579 -90 1583 -88
rect 1579 -92 1580 -90
rect 1582 -92 1583 -90
rect 1569 -99 1573 -98
rect 1569 -101 1570 -99
rect 1572 -101 1573 -99
rect 1521 -103 1561 -102
rect 1569 -103 1573 -101
rect 1579 -102 1583 -92
rect 1612 -78 1630 -77
rect 1612 -80 1614 -78
rect 1616 -80 1630 -78
rect 1612 -81 1630 -80
rect 1626 -87 1630 -81
rect 1626 -89 1627 -87
rect 1629 -89 1630 -87
rect 1605 -94 1611 -93
rect 1521 -105 1535 -103
rect 1537 -105 1561 -103
rect 1521 -106 1561 -105
rect 1577 -106 1583 -102
rect 1534 -110 1538 -106
rect 1557 -110 1581 -106
rect 1626 -102 1630 -89
rect 1615 -106 1630 -102
rect 1615 -110 1619 -106
rect 1633 -110 1634 -99
rect 1666 -78 1670 -74
rect 1681 -77 1682 -75
rect 1666 -82 1678 -78
rect 1674 -87 1678 -82
rect 1674 -89 1675 -87
rect 1677 -89 1678 -87
rect 1674 -101 1678 -89
rect 1661 -104 1678 -101
rect 1661 -106 1662 -104
rect 1664 -105 1678 -104
rect 1664 -106 1665 -105
rect 1403 -120 1409 -111
rect 1469 -111 1475 -110
rect 1469 -113 1471 -111
rect 1473 -113 1475 -111
rect 1434 -118 1440 -117
rect 1434 -120 1436 -118
rect 1438 -120 1440 -118
rect 1469 -118 1475 -113
rect 1482 -112 1483 -110
rect 1485 -112 1486 -110
rect 1482 -114 1486 -112
rect 1491 -111 1497 -110
rect 1491 -113 1493 -111
rect 1495 -113 1497 -111
rect 1469 -120 1471 -118
rect 1473 -120 1475 -118
rect 1491 -118 1497 -113
rect 1491 -120 1493 -118
rect 1495 -120 1497 -118
rect 1523 -111 1529 -110
rect 1523 -113 1525 -111
rect 1527 -113 1529 -111
rect 1523 -118 1529 -113
rect 1534 -112 1535 -110
rect 1537 -112 1538 -110
rect 1534 -114 1538 -112
rect 1545 -111 1551 -110
rect 1545 -113 1547 -111
rect 1549 -113 1551 -111
rect 1523 -120 1525 -118
rect 1527 -120 1529 -118
rect 1545 -118 1551 -113
rect 1602 -111 1619 -110
rect 1602 -113 1604 -111
rect 1606 -113 1619 -111
rect 1602 -114 1619 -113
rect 1650 -111 1656 -110
rect 1650 -113 1652 -111
rect 1654 -113 1656 -111
rect 1545 -120 1547 -118
rect 1549 -120 1551 -118
rect 1580 -118 1586 -117
rect 1580 -120 1582 -118
rect 1584 -120 1586 -118
rect 1621 -118 1627 -117
rect 1621 -120 1623 -118
rect 1625 -120 1627 -118
rect 1650 -120 1656 -113
rect 1661 -111 1665 -106
rect 1701 -71 1705 -69
rect 1710 -70 1735 -69
rect 1819 -70 1844 -69
rect 1710 -72 1712 -70
rect 1714 -71 1735 -70
rect 1714 -72 1732 -71
rect 1710 -73 1732 -72
rect 1734 -73 1735 -71
rect 1711 -78 1726 -77
rect 1711 -79 1722 -78
rect 1697 -80 1722 -79
rect 1724 -80 1726 -78
rect 1697 -82 1699 -80
rect 1701 -81 1726 -80
rect 1731 -78 1735 -73
rect 1740 -71 1750 -70
rect 1740 -73 1742 -71
rect 1744 -73 1750 -71
rect 1740 -74 1750 -73
rect 1731 -80 1732 -78
rect 1734 -80 1735 -78
rect 1701 -82 1715 -81
rect 1731 -82 1735 -80
rect 1697 -83 1715 -82
rect 1704 -90 1708 -88
rect 1704 -92 1705 -90
rect 1707 -92 1708 -90
rect 1704 -102 1708 -92
rect 1711 -94 1715 -83
rect 1746 -78 1750 -74
rect 1746 -82 1766 -78
rect 1762 -85 1766 -82
rect 1754 -87 1758 -85
rect 1754 -89 1755 -87
rect 1757 -89 1758 -87
rect 1754 -94 1758 -89
rect 1762 -87 1768 -85
rect 1762 -89 1765 -87
rect 1767 -89 1768 -87
rect 1762 -91 1768 -89
rect 1711 -98 1718 -94
rect 1714 -99 1718 -98
rect 1714 -101 1715 -99
rect 1717 -101 1718 -99
rect 1704 -106 1710 -102
rect 1714 -103 1718 -101
rect 1762 -102 1766 -91
rect 1726 -103 1766 -102
rect 1726 -105 1750 -103
rect 1752 -105 1766 -103
rect 1726 -106 1766 -105
rect 1661 -113 1662 -111
rect 1664 -113 1665 -111
rect 1661 -115 1665 -113
rect 1670 -109 1676 -108
rect 1670 -111 1672 -109
rect 1674 -111 1676 -109
rect 1706 -110 1730 -106
rect 1749 -110 1753 -106
rect 1804 -71 1814 -70
rect 1804 -73 1810 -71
rect 1812 -73 1814 -71
rect 1804 -74 1814 -73
rect 1819 -71 1840 -70
rect 1819 -73 1820 -71
rect 1822 -72 1840 -71
rect 1842 -72 1844 -70
rect 1849 -71 1853 -69
rect 1822 -73 1844 -72
rect 1926 -70 1932 -64
rect 1987 -67 1991 -64
rect 2043 -66 2045 -64
rect 2047 -66 2049 -64
rect 2043 -67 2049 -66
rect 2077 -66 2079 -64
rect 2081 -66 2083 -64
rect 2077 -67 2083 -66
rect 2135 -67 2139 -64
rect 1987 -69 1988 -67
rect 1990 -69 1991 -67
rect 2135 -69 2136 -67
rect 2138 -69 2139 -67
rect 2155 -65 2161 -64
rect 2155 -67 2157 -65
rect 2159 -67 2161 -65
rect 2155 -68 2161 -67
rect 2174 -65 2180 -64
rect 2174 -67 2176 -65
rect 2178 -67 2180 -65
rect 2174 -68 2180 -67
rect 1926 -72 1928 -70
rect 1930 -72 1932 -70
rect 1926 -73 1932 -72
rect 1939 -73 1943 -71
rect 1804 -78 1808 -74
rect 1788 -82 1808 -78
rect 1788 -85 1792 -82
rect 1786 -87 1792 -85
rect 1786 -89 1787 -87
rect 1789 -89 1792 -87
rect 1786 -91 1792 -89
rect 1788 -102 1792 -91
rect 1796 -87 1800 -85
rect 1819 -78 1823 -73
rect 1939 -75 1940 -73
rect 1942 -75 1943 -73
rect 1819 -80 1820 -78
rect 1822 -80 1823 -78
rect 1819 -82 1823 -80
rect 1828 -78 1843 -77
rect 1828 -80 1830 -78
rect 1832 -79 1843 -78
rect 1832 -80 1857 -79
rect 1828 -81 1853 -80
rect 1839 -82 1853 -81
rect 1855 -82 1857 -80
rect 1839 -83 1857 -82
rect 1796 -89 1797 -87
rect 1799 -89 1800 -87
rect 1796 -94 1800 -89
rect 1839 -94 1843 -83
rect 1836 -98 1843 -94
rect 1846 -90 1850 -88
rect 1846 -92 1847 -90
rect 1849 -92 1850 -90
rect 1836 -99 1840 -98
rect 1836 -101 1837 -99
rect 1839 -101 1840 -99
rect 1788 -103 1828 -102
rect 1836 -103 1840 -101
rect 1846 -102 1850 -92
rect 1879 -78 1897 -77
rect 1879 -80 1881 -78
rect 1883 -80 1897 -78
rect 1879 -81 1897 -80
rect 1893 -87 1897 -81
rect 1893 -89 1894 -87
rect 1896 -89 1897 -87
rect 1872 -94 1878 -93
rect 1788 -105 1802 -103
rect 1804 -105 1828 -103
rect 1788 -106 1828 -105
rect 1844 -106 1850 -102
rect 1801 -110 1805 -106
rect 1824 -110 1848 -106
rect 1893 -102 1897 -89
rect 1882 -106 1897 -102
rect 1882 -110 1886 -106
rect 1900 -110 1901 -99
rect 1913 -78 1917 -76
rect 1913 -80 1914 -78
rect 1916 -80 1917 -78
rect 1913 -86 1917 -80
rect 1939 -78 1943 -75
rect 1939 -82 1963 -78
rect 1913 -90 1924 -86
rect 1670 -120 1676 -111
rect 1736 -111 1742 -110
rect 1736 -113 1738 -111
rect 1740 -113 1742 -111
rect 1701 -118 1707 -117
rect 1701 -120 1703 -118
rect 1705 -120 1707 -118
rect 1736 -118 1742 -113
rect 1749 -112 1750 -110
rect 1752 -112 1753 -110
rect 1749 -114 1753 -112
rect 1758 -111 1764 -110
rect 1758 -113 1760 -111
rect 1762 -113 1764 -111
rect 1736 -120 1738 -118
rect 1740 -120 1742 -118
rect 1758 -118 1764 -113
rect 1758 -120 1760 -118
rect 1762 -120 1764 -118
rect 1790 -111 1796 -110
rect 1790 -113 1792 -111
rect 1794 -113 1796 -111
rect 1790 -118 1796 -113
rect 1801 -112 1802 -110
rect 1804 -112 1805 -110
rect 1801 -114 1805 -112
rect 1812 -111 1818 -110
rect 1812 -113 1814 -111
rect 1816 -113 1818 -111
rect 1790 -120 1792 -118
rect 1794 -120 1796 -118
rect 1812 -118 1818 -113
rect 1869 -111 1886 -110
rect 1869 -113 1871 -111
rect 1873 -113 1886 -111
rect 1869 -114 1886 -113
rect 1920 -96 1924 -90
rect 1959 -86 1963 -82
rect 1939 -87 1955 -86
rect 1939 -89 1951 -87
rect 1953 -89 1955 -87
rect 1939 -90 1955 -89
rect 1959 -88 1964 -86
rect 1959 -90 1961 -88
rect 1963 -90 1964 -88
rect 1939 -96 1943 -90
rect 1959 -92 1964 -90
rect 1959 -94 1963 -92
rect 1920 -97 1943 -96
rect 1920 -99 1922 -97
rect 1924 -99 1943 -97
rect 1920 -100 1943 -99
rect 1931 -111 1935 -109
rect 1931 -113 1932 -111
rect 1934 -113 1935 -111
rect 1812 -120 1814 -118
rect 1816 -120 1818 -118
rect 1847 -118 1853 -117
rect 1847 -120 1849 -118
rect 1851 -120 1853 -118
rect 1888 -118 1894 -117
rect 1888 -120 1890 -118
rect 1892 -120 1894 -118
rect 1931 -118 1935 -113
rect 1939 -111 1943 -100
rect 1947 -97 1963 -94
rect 1947 -99 1948 -97
rect 1950 -98 1963 -97
rect 1950 -99 1951 -98
rect 1947 -104 1951 -99
rect 1947 -106 1948 -104
rect 1950 -106 1951 -104
rect 1947 -108 1951 -106
rect 1987 -71 1991 -69
rect 1996 -70 2021 -69
rect 2105 -70 2130 -69
rect 1996 -72 1998 -70
rect 2000 -71 2021 -70
rect 2000 -72 2018 -71
rect 1996 -73 2018 -72
rect 2020 -73 2021 -71
rect 1997 -78 2012 -77
rect 1997 -79 2008 -78
rect 1983 -80 2008 -79
rect 2010 -80 2012 -78
rect 1983 -82 1985 -80
rect 1987 -81 2012 -80
rect 2017 -78 2021 -73
rect 2026 -71 2036 -70
rect 2026 -73 2028 -71
rect 2030 -73 2036 -71
rect 2026 -74 2036 -73
rect 2017 -80 2018 -78
rect 2020 -80 2021 -78
rect 1987 -82 2001 -81
rect 2017 -82 2021 -80
rect 1983 -83 2001 -82
rect 1990 -90 1994 -88
rect 1990 -92 1991 -90
rect 1993 -92 1994 -90
rect 1990 -102 1994 -92
rect 1997 -94 2001 -83
rect 2032 -78 2036 -74
rect 2032 -82 2052 -78
rect 2048 -85 2052 -82
rect 2040 -87 2044 -85
rect 2040 -89 2041 -87
rect 2043 -89 2044 -87
rect 2040 -94 2044 -89
rect 2048 -87 2054 -85
rect 2048 -89 2051 -87
rect 2053 -89 2054 -87
rect 2048 -91 2054 -89
rect 1997 -98 2004 -94
rect 2000 -99 2004 -98
rect 2000 -101 2001 -99
rect 2003 -101 2004 -99
rect 1990 -106 1996 -102
rect 2000 -103 2004 -101
rect 2048 -102 2052 -91
rect 2012 -103 2052 -102
rect 2012 -105 2036 -103
rect 2038 -105 2052 -103
rect 2012 -106 2052 -105
rect 1992 -110 2016 -106
rect 2035 -110 2039 -106
rect 2090 -71 2100 -70
rect 2090 -73 2096 -71
rect 2098 -73 2100 -71
rect 2090 -74 2100 -73
rect 2105 -71 2126 -70
rect 2105 -73 2106 -71
rect 2108 -72 2126 -71
rect 2128 -72 2130 -70
rect 2135 -71 2139 -69
rect 2108 -73 2130 -72
rect 2199 -72 2205 -71
rect 2090 -78 2094 -74
rect 2074 -82 2094 -78
rect 2074 -85 2078 -82
rect 2072 -87 2078 -85
rect 2072 -89 2073 -87
rect 2075 -89 2078 -87
rect 2072 -91 2078 -89
rect 2074 -102 2078 -91
rect 2082 -87 2086 -85
rect 2105 -78 2109 -73
rect 2105 -80 2106 -78
rect 2108 -80 2109 -78
rect 2105 -82 2109 -80
rect 2114 -78 2129 -77
rect 2114 -80 2116 -78
rect 2118 -79 2129 -78
rect 2118 -80 2143 -79
rect 2114 -81 2139 -80
rect 2125 -82 2139 -81
rect 2141 -82 2143 -80
rect 2125 -83 2143 -82
rect 2082 -89 2083 -87
rect 2085 -89 2086 -87
rect 2082 -94 2086 -89
rect 2125 -94 2129 -83
rect 2122 -98 2129 -94
rect 2132 -90 2136 -88
rect 2132 -92 2133 -90
rect 2135 -92 2136 -90
rect 2122 -99 2126 -98
rect 2122 -101 2123 -99
rect 2125 -101 2126 -99
rect 2074 -103 2114 -102
rect 2122 -103 2126 -101
rect 2132 -102 2136 -92
rect 2199 -74 2201 -72
rect 2203 -74 2205 -72
rect 2199 -75 2205 -74
rect 2209 -72 2215 -64
rect 2209 -74 2211 -72
rect 2213 -74 2215 -72
rect 2226 -70 2241 -69
rect 2226 -72 2228 -70
rect 2230 -72 2241 -70
rect 2226 -73 2241 -72
rect 2209 -75 2215 -74
rect 2165 -78 2183 -77
rect 2165 -80 2167 -78
rect 2169 -80 2183 -78
rect 2165 -81 2183 -80
rect 2179 -87 2183 -81
rect 2179 -89 2180 -87
rect 2182 -89 2183 -87
rect 2158 -94 2164 -93
rect 2074 -105 2088 -103
rect 2090 -105 2114 -103
rect 2074 -106 2114 -105
rect 2130 -106 2136 -102
rect 2087 -110 2091 -106
rect 2110 -110 2134 -106
rect 2179 -102 2183 -89
rect 2168 -106 2183 -102
rect 2168 -110 2172 -106
rect 2186 -110 2187 -99
rect 2199 -95 2203 -75
rect 2237 -78 2241 -73
rect 2244 -70 2248 -64
rect 2244 -72 2245 -70
rect 2247 -72 2248 -70
rect 2244 -74 2248 -72
rect 2223 -81 2234 -79
rect 2223 -83 2231 -81
rect 2233 -83 2234 -81
rect 2237 -80 2251 -78
rect 2237 -82 2252 -80
rect 2223 -85 2234 -83
rect 2247 -84 2249 -82
rect 2251 -84 2252 -82
rect 2223 -95 2227 -85
rect 2247 -86 2252 -84
rect 2199 -96 2227 -95
rect 2199 -98 2201 -96
rect 2203 -97 2227 -96
rect 2203 -98 2224 -97
rect 2199 -99 2224 -98
rect 2226 -99 2227 -97
rect 2243 -96 2244 -90
rect 2223 -101 2227 -99
rect 2022 -111 2028 -110
rect 1939 -112 1972 -111
rect 1939 -114 1968 -112
rect 1970 -114 1972 -112
rect 1939 -115 1972 -114
rect 2022 -113 2024 -111
rect 2026 -113 2028 -111
rect 1931 -120 1932 -118
rect 1934 -120 1935 -118
rect 1987 -118 1993 -117
rect 1987 -120 1989 -118
rect 1991 -120 1993 -118
rect 2022 -118 2028 -113
rect 2035 -112 2036 -110
rect 2038 -112 2039 -110
rect 2035 -114 2039 -112
rect 2044 -111 2050 -110
rect 2044 -113 2046 -111
rect 2048 -113 2050 -111
rect 2022 -120 2024 -118
rect 2026 -120 2028 -118
rect 2044 -118 2050 -113
rect 2044 -120 2046 -118
rect 2048 -120 2050 -118
rect 2076 -111 2082 -110
rect 2076 -113 2078 -111
rect 2080 -113 2082 -111
rect 2076 -118 2082 -113
rect 2087 -112 2088 -110
rect 2090 -112 2091 -110
rect 2087 -114 2091 -112
rect 2098 -111 2104 -110
rect 2098 -113 2100 -111
rect 2102 -113 2104 -111
rect 2076 -120 2078 -118
rect 2080 -120 2082 -118
rect 2098 -118 2104 -113
rect 2155 -111 2172 -110
rect 2155 -113 2157 -111
rect 2159 -113 2172 -111
rect 2155 -114 2172 -113
rect 2247 -103 2251 -86
rect 2235 -107 2251 -103
rect 2226 -108 2239 -107
rect 2226 -110 2228 -108
rect 2230 -110 2239 -108
rect 2267 -72 2273 -71
rect 2267 -74 2269 -72
rect 2271 -74 2273 -72
rect 2267 -75 2273 -74
rect 2277 -72 2283 -64
rect 2277 -74 2279 -72
rect 2281 -74 2283 -72
rect 2294 -70 2309 -69
rect 2294 -72 2296 -70
rect 2298 -72 2309 -70
rect 2294 -73 2309 -72
rect 2277 -75 2283 -74
rect 2267 -95 2271 -75
rect 2305 -78 2309 -73
rect 2312 -70 2316 -64
rect 2312 -72 2313 -70
rect 2315 -72 2316 -70
rect 2312 -74 2316 -72
rect 2291 -81 2302 -79
rect 2291 -83 2299 -81
rect 2301 -83 2302 -81
rect 2305 -80 2319 -78
rect 2305 -82 2320 -80
rect 2291 -85 2302 -83
rect 2315 -84 2317 -82
rect 2319 -84 2320 -82
rect 2291 -95 2295 -85
rect 2315 -86 2320 -84
rect 2267 -96 2295 -95
rect 2267 -98 2269 -96
rect 2271 -97 2295 -96
rect 2271 -98 2292 -97
rect 2267 -99 2292 -98
rect 2294 -99 2295 -97
rect 2311 -96 2312 -90
rect 2291 -101 2295 -99
rect 2226 -111 2239 -110
rect 2315 -103 2319 -86
rect 2303 -107 2319 -103
rect 2294 -108 2307 -107
rect 2294 -110 2296 -108
rect 2298 -110 2307 -108
rect 2294 -111 2307 -110
rect 2098 -120 2100 -118
rect 2102 -120 2104 -118
rect 2133 -118 2139 -117
rect 2133 -120 2135 -118
rect 2137 -120 2139 -118
rect 2174 -118 2180 -117
rect 2174 -120 2176 -118
rect 2178 -120 2180 -118
rect 2210 -118 2214 -116
rect 2210 -120 2211 -118
rect 2213 -120 2214 -118
rect 2243 -118 2249 -117
rect 2243 -120 2245 -118
rect 2247 -120 2249 -118
rect 2278 -118 2282 -116
rect 2278 -120 2279 -118
rect 2281 -120 2282 -118
rect 2311 -118 2317 -117
rect 2311 -120 2313 -118
rect 2315 -120 2317 -118
rect 8 -143 14 -136
rect 8 -145 10 -143
rect 12 -145 14 -143
rect 8 -146 14 -145
rect 19 -143 23 -141
rect 19 -145 20 -143
rect 22 -145 23 -143
rect 19 -150 23 -145
rect 28 -145 34 -136
rect 48 -143 54 -136
rect 48 -145 50 -143
rect 52 -145 54 -143
rect 28 -147 30 -145
rect 32 -147 34 -145
rect 28 -148 34 -147
rect 48 -146 54 -145
rect 59 -143 63 -141
rect 59 -145 60 -143
rect 62 -145 63 -143
rect 19 -152 20 -150
rect 22 -151 23 -150
rect 22 -152 36 -151
rect 19 -155 36 -152
rect 32 -167 36 -155
rect 59 -150 63 -145
rect 68 -145 74 -136
rect 99 -138 101 -136
rect 103 -138 105 -136
rect 99 -139 105 -138
rect 134 -138 136 -136
rect 138 -138 140 -136
rect 68 -147 70 -145
rect 72 -147 74 -145
rect 134 -143 140 -138
rect 156 -138 158 -136
rect 160 -138 162 -136
rect 134 -145 136 -143
rect 138 -145 140 -143
rect 134 -146 140 -145
rect 147 -144 151 -142
rect 147 -146 148 -144
rect 150 -146 151 -144
rect 156 -143 162 -138
rect 156 -145 158 -143
rect 160 -145 162 -143
rect 156 -146 162 -145
rect 188 -138 190 -136
rect 192 -138 194 -136
rect 188 -143 194 -138
rect 210 -138 212 -136
rect 214 -138 216 -136
rect 188 -145 190 -143
rect 192 -145 194 -143
rect 188 -146 194 -145
rect 199 -144 203 -142
rect 199 -146 200 -144
rect 202 -146 203 -144
rect 210 -143 216 -138
rect 245 -138 247 -136
rect 249 -138 251 -136
rect 245 -139 251 -138
rect 286 -138 288 -136
rect 290 -138 292 -136
rect 286 -139 292 -138
rect 210 -145 212 -143
rect 214 -145 216 -143
rect 210 -146 216 -145
rect 267 -143 284 -142
rect 267 -145 269 -143
rect 271 -145 284 -143
rect 267 -146 284 -145
rect 315 -143 321 -136
rect 315 -145 317 -143
rect 319 -145 321 -143
rect 315 -146 321 -145
rect 326 -143 330 -141
rect 326 -145 327 -143
rect 329 -145 330 -143
rect 68 -148 74 -147
rect 59 -152 60 -150
rect 62 -151 63 -150
rect 62 -152 76 -151
rect 59 -155 76 -152
rect 32 -169 33 -167
rect 35 -169 36 -167
rect 32 -174 36 -169
rect 24 -178 36 -174
rect 24 -182 28 -178
rect 39 -181 40 -179
rect 72 -167 76 -155
rect 72 -169 73 -167
rect 75 -169 76 -167
rect 72 -174 76 -169
rect 64 -178 76 -174
rect 8 -183 28 -182
rect 8 -185 10 -183
rect 12 -185 28 -183
rect 8 -186 28 -185
rect 64 -182 68 -178
rect 79 -181 80 -179
rect 48 -183 68 -182
rect 48 -185 50 -183
rect 52 -185 68 -183
rect 48 -186 68 -185
rect 104 -150 128 -146
rect 147 -150 151 -146
rect 102 -154 108 -150
rect 124 -151 164 -150
rect 124 -153 148 -151
rect 150 -153 164 -151
rect 102 -164 106 -154
rect 112 -155 116 -153
rect 124 -154 164 -153
rect 112 -157 113 -155
rect 115 -157 116 -155
rect 112 -158 116 -157
rect 102 -166 103 -164
rect 105 -166 106 -164
rect 102 -168 106 -166
rect 109 -162 116 -158
rect 109 -173 113 -162
rect 152 -167 156 -162
rect 152 -169 153 -167
rect 155 -169 156 -167
rect 95 -174 113 -173
rect 95 -176 97 -174
rect 99 -175 113 -174
rect 99 -176 124 -175
rect 95 -177 120 -176
rect 109 -178 120 -177
rect 122 -178 124 -176
rect 109 -179 124 -178
rect 129 -176 133 -174
rect 129 -178 130 -176
rect 132 -178 133 -176
rect 129 -183 133 -178
rect 152 -171 156 -169
rect 160 -165 164 -154
rect 160 -167 166 -165
rect 160 -169 163 -167
rect 165 -169 166 -167
rect 160 -171 166 -169
rect 160 -174 164 -171
rect 144 -178 164 -174
rect 144 -182 148 -178
rect 108 -184 130 -183
rect 99 -187 103 -185
rect 108 -186 110 -184
rect 112 -185 130 -184
rect 132 -185 133 -183
rect 112 -186 133 -185
rect 138 -183 148 -182
rect 138 -185 140 -183
rect 142 -185 148 -183
rect 138 -186 148 -185
rect 199 -150 203 -146
rect 222 -150 246 -146
rect 186 -151 226 -150
rect 186 -153 200 -151
rect 202 -153 226 -151
rect 186 -154 226 -153
rect 186 -165 190 -154
rect 234 -155 238 -153
rect 242 -154 248 -150
rect 234 -157 235 -155
rect 237 -157 238 -155
rect 234 -158 238 -157
rect 234 -162 241 -158
rect 184 -167 190 -165
rect 184 -169 185 -167
rect 187 -169 190 -167
rect 184 -171 190 -169
rect 194 -167 198 -162
rect 194 -169 195 -167
rect 197 -169 198 -167
rect 194 -171 198 -169
rect 186 -174 190 -171
rect 186 -178 206 -174
rect 202 -182 206 -178
rect 237 -173 241 -162
rect 244 -164 248 -154
rect 244 -166 245 -164
rect 247 -166 248 -164
rect 244 -168 248 -166
rect 237 -174 255 -173
rect 217 -176 221 -174
rect 237 -175 251 -174
rect 217 -178 218 -176
rect 220 -178 221 -176
rect 202 -183 212 -182
rect 202 -185 208 -183
rect 210 -185 212 -183
rect 202 -186 212 -185
rect 217 -183 221 -178
rect 226 -176 251 -175
rect 253 -176 255 -174
rect 226 -178 228 -176
rect 230 -177 255 -176
rect 230 -178 241 -177
rect 226 -179 241 -178
rect 280 -150 284 -146
rect 280 -154 295 -150
rect 270 -163 276 -162
rect 291 -167 295 -154
rect 298 -157 299 -146
rect 291 -169 292 -167
rect 294 -169 295 -167
rect 291 -175 295 -169
rect 326 -150 330 -145
rect 335 -145 341 -136
rect 366 -138 368 -136
rect 370 -138 372 -136
rect 366 -139 372 -138
rect 401 -138 403 -136
rect 405 -138 407 -136
rect 335 -147 337 -145
rect 339 -147 341 -145
rect 401 -143 407 -138
rect 423 -138 425 -136
rect 427 -138 429 -136
rect 401 -145 403 -143
rect 405 -145 407 -143
rect 401 -146 407 -145
rect 414 -144 418 -142
rect 414 -146 415 -144
rect 417 -146 418 -144
rect 423 -143 429 -138
rect 423 -145 425 -143
rect 427 -145 429 -143
rect 423 -146 429 -145
rect 455 -138 457 -136
rect 459 -138 461 -136
rect 455 -143 461 -138
rect 477 -138 479 -136
rect 481 -138 483 -136
rect 455 -145 457 -143
rect 459 -145 461 -143
rect 455 -146 461 -145
rect 466 -144 470 -142
rect 466 -146 467 -144
rect 469 -146 470 -144
rect 477 -143 483 -138
rect 512 -138 514 -136
rect 516 -138 518 -136
rect 512 -139 518 -138
rect 553 -138 555 -136
rect 557 -138 559 -136
rect 553 -139 559 -138
rect 477 -145 479 -143
rect 481 -145 483 -143
rect 477 -146 483 -145
rect 534 -143 551 -142
rect 534 -145 536 -143
rect 538 -145 551 -143
rect 534 -146 551 -145
rect 582 -143 588 -136
rect 582 -145 584 -143
rect 586 -145 588 -143
rect 582 -146 588 -145
rect 593 -143 597 -141
rect 593 -145 594 -143
rect 596 -145 597 -143
rect 335 -148 341 -147
rect 326 -152 327 -150
rect 329 -151 330 -150
rect 329 -152 343 -151
rect 326 -155 343 -152
rect 277 -176 295 -175
rect 277 -178 279 -176
rect 281 -178 295 -176
rect 277 -179 295 -178
rect 339 -167 343 -155
rect 339 -169 340 -167
rect 342 -169 343 -167
rect 339 -174 343 -169
rect 331 -178 343 -174
rect 331 -182 335 -178
rect 346 -181 347 -179
rect 217 -185 218 -183
rect 220 -184 242 -183
rect 220 -185 238 -184
rect 217 -186 238 -185
rect 240 -186 242 -184
rect 108 -187 133 -186
rect 217 -187 242 -186
rect 247 -187 251 -185
rect 315 -183 335 -182
rect 315 -185 317 -183
rect 319 -185 335 -183
rect 315 -186 335 -185
rect 371 -150 395 -146
rect 414 -150 418 -146
rect 369 -154 375 -150
rect 391 -151 431 -150
rect 391 -153 415 -151
rect 417 -153 431 -151
rect 369 -164 373 -154
rect 379 -155 383 -153
rect 391 -154 431 -153
rect 379 -157 380 -155
rect 382 -157 383 -155
rect 379 -158 383 -157
rect 369 -166 370 -164
rect 372 -166 373 -164
rect 369 -168 373 -166
rect 376 -162 383 -158
rect 376 -173 380 -162
rect 419 -167 423 -162
rect 419 -169 420 -167
rect 422 -169 423 -167
rect 362 -174 380 -173
rect 362 -176 364 -174
rect 366 -175 380 -174
rect 366 -176 391 -175
rect 362 -177 387 -176
rect 376 -178 387 -177
rect 389 -178 391 -176
rect 376 -179 391 -178
rect 396 -176 400 -174
rect 396 -178 397 -176
rect 399 -178 400 -176
rect 396 -183 400 -178
rect 419 -171 423 -169
rect 427 -165 431 -154
rect 427 -167 433 -165
rect 427 -169 430 -167
rect 432 -169 433 -167
rect 427 -171 433 -169
rect 427 -174 431 -171
rect 411 -178 431 -174
rect 411 -182 415 -178
rect 375 -184 397 -183
rect 366 -187 370 -185
rect 375 -186 377 -184
rect 379 -185 397 -184
rect 399 -185 400 -183
rect 379 -186 400 -185
rect 405 -183 415 -182
rect 405 -185 407 -183
rect 409 -185 415 -183
rect 405 -186 415 -185
rect 466 -150 470 -146
rect 489 -150 513 -146
rect 453 -151 493 -150
rect 453 -153 467 -151
rect 469 -153 493 -151
rect 453 -154 493 -153
rect 453 -165 457 -154
rect 501 -155 505 -153
rect 509 -154 515 -150
rect 501 -157 502 -155
rect 504 -157 505 -155
rect 501 -158 505 -157
rect 501 -162 508 -158
rect 451 -167 457 -165
rect 451 -169 452 -167
rect 454 -169 457 -167
rect 451 -171 457 -169
rect 461 -167 465 -162
rect 461 -169 462 -167
rect 464 -169 465 -167
rect 461 -171 465 -169
rect 453 -174 457 -171
rect 453 -178 473 -174
rect 469 -182 473 -178
rect 504 -173 508 -162
rect 511 -164 515 -154
rect 511 -166 512 -164
rect 514 -166 515 -164
rect 511 -168 515 -166
rect 504 -174 522 -173
rect 484 -176 488 -174
rect 504 -175 518 -174
rect 484 -178 485 -176
rect 487 -178 488 -176
rect 469 -183 479 -182
rect 469 -185 475 -183
rect 477 -185 479 -183
rect 469 -186 479 -185
rect 484 -183 488 -178
rect 493 -176 518 -175
rect 520 -176 522 -174
rect 493 -178 495 -176
rect 497 -177 522 -176
rect 497 -178 508 -177
rect 493 -179 508 -178
rect 547 -150 551 -146
rect 547 -154 562 -150
rect 537 -163 543 -162
rect 558 -167 562 -154
rect 565 -157 566 -146
rect 558 -169 559 -167
rect 561 -169 562 -167
rect 558 -175 562 -169
rect 593 -150 597 -145
rect 602 -145 608 -136
rect 633 -138 635 -136
rect 637 -138 639 -136
rect 633 -139 639 -138
rect 668 -138 670 -136
rect 672 -138 674 -136
rect 602 -147 604 -145
rect 606 -147 608 -145
rect 668 -143 674 -138
rect 690 -138 692 -136
rect 694 -138 696 -136
rect 668 -145 670 -143
rect 672 -145 674 -143
rect 668 -146 674 -145
rect 681 -144 685 -142
rect 681 -146 682 -144
rect 684 -146 685 -144
rect 690 -143 696 -138
rect 690 -145 692 -143
rect 694 -145 696 -143
rect 690 -146 696 -145
rect 722 -138 724 -136
rect 726 -138 728 -136
rect 722 -143 728 -138
rect 744 -138 746 -136
rect 748 -138 750 -136
rect 722 -145 724 -143
rect 726 -145 728 -143
rect 722 -146 728 -145
rect 733 -144 737 -142
rect 733 -146 734 -144
rect 736 -146 737 -144
rect 744 -143 750 -138
rect 779 -138 781 -136
rect 783 -138 785 -136
rect 779 -139 785 -138
rect 820 -138 822 -136
rect 824 -138 826 -136
rect 820 -139 826 -138
rect 744 -145 746 -143
rect 748 -145 750 -143
rect 744 -146 750 -145
rect 801 -143 818 -142
rect 801 -145 803 -143
rect 805 -145 818 -143
rect 801 -146 818 -145
rect 849 -143 855 -136
rect 849 -145 851 -143
rect 853 -145 855 -143
rect 849 -146 855 -145
rect 860 -143 864 -141
rect 860 -145 861 -143
rect 863 -145 864 -143
rect 602 -148 608 -147
rect 593 -152 594 -150
rect 596 -151 597 -150
rect 596 -152 610 -151
rect 593 -155 610 -152
rect 544 -176 562 -175
rect 544 -178 546 -176
rect 548 -178 562 -176
rect 544 -179 562 -178
rect 606 -167 610 -155
rect 606 -169 607 -167
rect 609 -169 610 -167
rect 606 -174 610 -169
rect 598 -178 610 -174
rect 598 -182 602 -178
rect 613 -181 614 -179
rect 484 -185 485 -183
rect 487 -184 509 -183
rect 487 -185 505 -184
rect 484 -186 505 -185
rect 507 -186 509 -184
rect 375 -187 400 -186
rect 484 -187 509 -186
rect 514 -187 518 -185
rect 582 -183 602 -182
rect 582 -185 584 -183
rect 586 -185 602 -183
rect 582 -186 602 -185
rect 638 -150 662 -146
rect 681 -150 685 -146
rect 636 -154 642 -150
rect 658 -151 698 -150
rect 658 -153 682 -151
rect 684 -153 698 -151
rect 636 -164 640 -154
rect 646 -155 650 -153
rect 658 -154 698 -153
rect 646 -157 647 -155
rect 649 -157 650 -155
rect 646 -158 650 -157
rect 636 -166 637 -164
rect 639 -166 640 -164
rect 636 -168 640 -166
rect 643 -162 650 -158
rect 643 -173 647 -162
rect 686 -167 690 -162
rect 686 -169 687 -167
rect 689 -169 690 -167
rect 629 -174 647 -173
rect 629 -176 631 -174
rect 633 -175 647 -174
rect 633 -176 658 -175
rect 629 -177 654 -176
rect 643 -178 654 -177
rect 656 -178 658 -176
rect 643 -179 658 -178
rect 663 -176 667 -174
rect 663 -178 664 -176
rect 666 -178 667 -176
rect 663 -183 667 -178
rect 686 -171 690 -169
rect 694 -165 698 -154
rect 694 -167 700 -165
rect 694 -169 697 -167
rect 699 -169 700 -167
rect 694 -171 700 -169
rect 694 -174 698 -171
rect 678 -178 698 -174
rect 678 -182 682 -178
rect 642 -184 664 -183
rect 633 -187 637 -185
rect 642 -186 644 -184
rect 646 -185 664 -184
rect 666 -185 667 -183
rect 646 -186 667 -185
rect 672 -183 682 -182
rect 672 -185 674 -183
rect 676 -185 682 -183
rect 672 -186 682 -185
rect 733 -150 737 -146
rect 756 -150 780 -146
rect 720 -151 760 -150
rect 720 -153 734 -151
rect 736 -153 760 -151
rect 720 -154 760 -153
rect 720 -165 724 -154
rect 768 -155 772 -153
rect 776 -154 782 -150
rect 768 -157 769 -155
rect 771 -157 772 -155
rect 768 -158 772 -157
rect 768 -162 775 -158
rect 718 -167 724 -165
rect 718 -169 719 -167
rect 721 -169 724 -167
rect 718 -171 724 -169
rect 728 -167 732 -162
rect 728 -169 729 -167
rect 731 -169 732 -167
rect 728 -171 732 -169
rect 720 -174 724 -171
rect 720 -178 740 -174
rect 736 -182 740 -178
rect 771 -173 775 -162
rect 778 -164 782 -154
rect 778 -166 779 -164
rect 781 -166 782 -164
rect 778 -168 782 -166
rect 771 -174 789 -173
rect 751 -176 755 -174
rect 771 -175 785 -174
rect 751 -178 752 -176
rect 754 -178 755 -176
rect 736 -183 746 -182
rect 736 -185 742 -183
rect 744 -185 746 -183
rect 736 -186 746 -185
rect 751 -183 755 -178
rect 760 -176 785 -175
rect 787 -176 789 -174
rect 760 -178 762 -176
rect 764 -177 789 -176
rect 764 -178 775 -177
rect 760 -179 775 -178
rect 814 -150 818 -146
rect 814 -154 829 -150
rect 804 -163 810 -162
rect 825 -167 829 -154
rect 832 -157 833 -146
rect 825 -169 826 -167
rect 828 -169 829 -167
rect 825 -175 829 -169
rect 860 -150 864 -145
rect 869 -145 875 -136
rect 900 -138 902 -136
rect 904 -138 906 -136
rect 900 -139 906 -138
rect 935 -138 937 -136
rect 939 -138 941 -136
rect 869 -147 871 -145
rect 873 -147 875 -145
rect 935 -143 941 -138
rect 957 -138 959 -136
rect 961 -138 963 -136
rect 935 -145 937 -143
rect 939 -145 941 -143
rect 935 -146 941 -145
rect 948 -144 952 -142
rect 948 -146 949 -144
rect 951 -146 952 -144
rect 957 -143 963 -138
rect 957 -145 959 -143
rect 961 -145 963 -143
rect 957 -146 963 -145
rect 989 -138 991 -136
rect 993 -138 995 -136
rect 989 -143 995 -138
rect 1011 -138 1013 -136
rect 1015 -138 1017 -136
rect 989 -145 991 -143
rect 993 -145 995 -143
rect 989 -146 995 -145
rect 1000 -144 1004 -142
rect 1000 -146 1001 -144
rect 1003 -146 1004 -144
rect 1011 -143 1017 -138
rect 1046 -138 1048 -136
rect 1050 -138 1052 -136
rect 1046 -139 1052 -138
rect 1087 -138 1089 -136
rect 1091 -138 1093 -136
rect 1087 -139 1093 -138
rect 1011 -145 1013 -143
rect 1015 -145 1017 -143
rect 1011 -146 1017 -145
rect 1068 -143 1085 -142
rect 1068 -145 1070 -143
rect 1072 -145 1085 -143
rect 1068 -146 1085 -145
rect 1116 -143 1122 -136
rect 1116 -145 1118 -143
rect 1120 -145 1122 -143
rect 1116 -146 1122 -145
rect 1127 -143 1131 -141
rect 1127 -145 1128 -143
rect 1130 -145 1131 -143
rect 869 -148 875 -147
rect 860 -152 861 -150
rect 863 -151 864 -150
rect 863 -152 877 -151
rect 860 -155 877 -152
rect 811 -176 829 -175
rect 811 -178 813 -176
rect 815 -178 829 -176
rect 811 -179 829 -178
rect 873 -167 877 -155
rect 873 -169 874 -167
rect 876 -169 877 -167
rect 873 -174 877 -169
rect 865 -178 877 -174
rect 865 -182 869 -178
rect 880 -181 881 -179
rect 751 -185 752 -183
rect 754 -184 776 -183
rect 754 -185 772 -184
rect 751 -186 772 -185
rect 774 -186 776 -184
rect 642 -187 667 -186
rect 751 -187 776 -186
rect 781 -187 785 -185
rect 849 -183 869 -182
rect 849 -185 851 -183
rect 853 -185 869 -183
rect 849 -186 869 -185
rect 905 -150 929 -146
rect 948 -150 952 -146
rect 903 -154 909 -150
rect 925 -151 965 -150
rect 925 -153 949 -151
rect 951 -153 965 -151
rect 903 -164 907 -154
rect 913 -155 917 -153
rect 925 -154 965 -153
rect 913 -157 914 -155
rect 916 -157 917 -155
rect 913 -158 917 -157
rect 903 -166 904 -164
rect 906 -166 907 -164
rect 903 -168 907 -166
rect 910 -162 917 -158
rect 910 -173 914 -162
rect 953 -167 957 -162
rect 953 -169 954 -167
rect 956 -169 957 -167
rect 896 -174 914 -173
rect 896 -176 898 -174
rect 900 -175 914 -174
rect 900 -176 925 -175
rect 896 -177 921 -176
rect 910 -178 921 -177
rect 923 -178 925 -176
rect 910 -179 925 -178
rect 930 -176 934 -174
rect 930 -178 931 -176
rect 933 -178 934 -176
rect 930 -183 934 -178
rect 953 -171 957 -169
rect 961 -165 965 -154
rect 961 -167 967 -165
rect 961 -169 964 -167
rect 966 -169 967 -167
rect 961 -171 967 -169
rect 961 -174 965 -171
rect 945 -178 965 -174
rect 945 -182 949 -178
rect 909 -184 931 -183
rect 900 -187 904 -185
rect 909 -186 911 -184
rect 913 -185 931 -184
rect 933 -185 934 -183
rect 913 -186 934 -185
rect 939 -183 949 -182
rect 939 -185 941 -183
rect 943 -185 949 -183
rect 939 -186 949 -185
rect 1000 -150 1004 -146
rect 1023 -150 1047 -146
rect 987 -151 1027 -150
rect 987 -153 1001 -151
rect 1003 -153 1027 -151
rect 987 -154 1027 -153
rect 987 -165 991 -154
rect 1035 -155 1039 -153
rect 1043 -154 1049 -150
rect 1035 -157 1036 -155
rect 1038 -157 1039 -155
rect 1035 -158 1039 -157
rect 1035 -162 1042 -158
rect 985 -167 991 -165
rect 985 -169 986 -167
rect 988 -169 991 -167
rect 985 -171 991 -169
rect 995 -167 999 -162
rect 995 -169 996 -167
rect 998 -169 999 -167
rect 995 -171 999 -169
rect 987 -174 991 -171
rect 987 -178 1007 -174
rect 1003 -182 1007 -178
rect 1038 -173 1042 -162
rect 1045 -164 1049 -154
rect 1045 -166 1046 -164
rect 1048 -166 1049 -164
rect 1045 -168 1049 -166
rect 1038 -174 1056 -173
rect 1018 -176 1022 -174
rect 1038 -175 1052 -174
rect 1018 -178 1019 -176
rect 1021 -178 1022 -176
rect 1003 -183 1013 -182
rect 1003 -185 1009 -183
rect 1011 -185 1013 -183
rect 1003 -186 1013 -185
rect 1018 -183 1022 -178
rect 1027 -176 1052 -175
rect 1054 -176 1056 -174
rect 1027 -178 1029 -176
rect 1031 -177 1056 -176
rect 1031 -178 1042 -177
rect 1027 -179 1042 -178
rect 1081 -150 1085 -146
rect 1081 -154 1096 -150
rect 1071 -163 1077 -162
rect 1092 -167 1096 -154
rect 1099 -157 1100 -146
rect 1092 -169 1093 -167
rect 1095 -169 1096 -167
rect 1092 -175 1096 -169
rect 1127 -150 1131 -145
rect 1136 -145 1142 -136
rect 1167 -138 1169 -136
rect 1171 -138 1173 -136
rect 1167 -139 1173 -138
rect 1202 -138 1204 -136
rect 1206 -138 1208 -136
rect 1136 -147 1138 -145
rect 1140 -147 1142 -145
rect 1202 -143 1208 -138
rect 1224 -138 1226 -136
rect 1228 -138 1230 -136
rect 1202 -145 1204 -143
rect 1206 -145 1208 -143
rect 1202 -146 1208 -145
rect 1215 -144 1219 -142
rect 1215 -146 1216 -144
rect 1218 -146 1219 -144
rect 1224 -143 1230 -138
rect 1224 -145 1226 -143
rect 1228 -145 1230 -143
rect 1224 -146 1230 -145
rect 1256 -138 1258 -136
rect 1260 -138 1262 -136
rect 1256 -143 1262 -138
rect 1278 -138 1280 -136
rect 1282 -138 1284 -136
rect 1256 -145 1258 -143
rect 1260 -145 1262 -143
rect 1256 -146 1262 -145
rect 1267 -144 1271 -142
rect 1267 -146 1268 -144
rect 1270 -146 1271 -144
rect 1278 -143 1284 -138
rect 1313 -138 1315 -136
rect 1317 -138 1319 -136
rect 1313 -139 1319 -138
rect 1354 -138 1356 -136
rect 1358 -138 1360 -136
rect 1354 -139 1360 -138
rect 1278 -145 1280 -143
rect 1282 -145 1284 -143
rect 1278 -146 1284 -145
rect 1335 -143 1352 -142
rect 1335 -145 1337 -143
rect 1339 -145 1352 -143
rect 1335 -146 1352 -145
rect 1383 -143 1389 -136
rect 1383 -145 1385 -143
rect 1387 -145 1389 -143
rect 1383 -146 1389 -145
rect 1394 -143 1398 -141
rect 1394 -145 1395 -143
rect 1397 -145 1398 -143
rect 1136 -148 1142 -147
rect 1127 -152 1128 -150
rect 1130 -151 1131 -150
rect 1130 -152 1144 -151
rect 1127 -155 1144 -152
rect 1078 -176 1096 -175
rect 1078 -178 1080 -176
rect 1082 -178 1096 -176
rect 1078 -179 1096 -178
rect 1140 -167 1144 -155
rect 1140 -169 1141 -167
rect 1143 -169 1144 -167
rect 1140 -174 1144 -169
rect 1132 -178 1144 -174
rect 1132 -182 1136 -178
rect 1147 -181 1148 -179
rect 1018 -185 1019 -183
rect 1021 -184 1043 -183
rect 1021 -185 1039 -184
rect 1018 -186 1039 -185
rect 1041 -186 1043 -184
rect 909 -187 934 -186
rect 1018 -187 1043 -186
rect 1048 -187 1052 -185
rect 1116 -183 1136 -182
rect 1116 -185 1118 -183
rect 1120 -185 1136 -183
rect 1116 -186 1136 -185
rect 1172 -150 1196 -146
rect 1215 -150 1219 -146
rect 1170 -154 1176 -150
rect 1192 -151 1232 -150
rect 1192 -153 1216 -151
rect 1218 -153 1232 -151
rect 1170 -164 1174 -154
rect 1180 -155 1184 -153
rect 1192 -154 1232 -153
rect 1180 -157 1181 -155
rect 1183 -157 1184 -155
rect 1180 -158 1184 -157
rect 1170 -166 1171 -164
rect 1173 -166 1174 -164
rect 1170 -168 1174 -166
rect 1177 -162 1184 -158
rect 1177 -173 1181 -162
rect 1220 -167 1224 -162
rect 1220 -169 1221 -167
rect 1223 -169 1224 -167
rect 1163 -174 1181 -173
rect 1163 -176 1165 -174
rect 1167 -175 1181 -174
rect 1167 -176 1192 -175
rect 1163 -177 1188 -176
rect 1177 -178 1188 -177
rect 1190 -178 1192 -176
rect 1177 -179 1192 -178
rect 1197 -176 1201 -174
rect 1197 -178 1198 -176
rect 1200 -178 1201 -176
rect 1197 -183 1201 -178
rect 1220 -171 1224 -169
rect 1228 -165 1232 -154
rect 1228 -167 1234 -165
rect 1228 -169 1231 -167
rect 1233 -169 1234 -167
rect 1228 -171 1234 -169
rect 1228 -174 1232 -171
rect 1212 -178 1232 -174
rect 1212 -182 1216 -178
rect 1176 -184 1198 -183
rect 1167 -187 1171 -185
rect 1176 -186 1178 -184
rect 1180 -185 1198 -184
rect 1200 -185 1201 -183
rect 1180 -186 1201 -185
rect 1206 -183 1216 -182
rect 1206 -185 1208 -183
rect 1210 -185 1216 -183
rect 1206 -186 1216 -185
rect 1267 -150 1271 -146
rect 1290 -150 1314 -146
rect 1254 -151 1294 -150
rect 1254 -153 1268 -151
rect 1270 -153 1294 -151
rect 1254 -154 1294 -153
rect 1254 -165 1258 -154
rect 1302 -155 1306 -153
rect 1310 -154 1316 -150
rect 1302 -157 1303 -155
rect 1305 -157 1306 -155
rect 1302 -158 1306 -157
rect 1302 -162 1309 -158
rect 1252 -167 1258 -165
rect 1252 -169 1253 -167
rect 1255 -169 1258 -167
rect 1252 -171 1258 -169
rect 1262 -167 1266 -162
rect 1262 -169 1263 -167
rect 1265 -169 1266 -167
rect 1262 -171 1266 -169
rect 1254 -174 1258 -171
rect 1254 -178 1274 -174
rect 1270 -182 1274 -178
rect 1305 -173 1309 -162
rect 1312 -164 1316 -154
rect 1312 -166 1313 -164
rect 1315 -166 1316 -164
rect 1312 -168 1316 -166
rect 1305 -174 1323 -173
rect 1285 -176 1289 -174
rect 1305 -175 1319 -174
rect 1285 -178 1286 -176
rect 1288 -178 1289 -176
rect 1270 -183 1280 -182
rect 1270 -185 1276 -183
rect 1278 -185 1280 -183
rect 1270 -186 1280 -185
rect 1285 -183 1289 -178
rect 1294 -176 1319 -175
rect 1321 -176 1323 -174
rect 1294 -178 1296 -176
rect 1298 -177 1323 -176
rect 1298 -178 1309 -177
rect 1294 -179 1309 -178
rect 1348 -150 1352 -146
rect 1348 -154 1363 -150
rect 1338 -163 1344 -162
rect 1359 -167 1363 -154
rect 1366 -157 1367 -146
rect 1359 -169 1360 -167
rect 1362 -169 1363 -167
rect 1359 -175 1363 -169
rect 1394 -150 1398 -145
rect 1403 -145 1409 -136
rect 1434 -138 1436 -136
rect 1438 -138 1440 -136
rect 1434 -139 1440 -138
rect 1469 -138 1471 -136
rect 1473 -138 1475 -136
rect 1403 -147 1405 -145
rect 1407 -147 1409 -145
rect 1469 -143 1475 -138
rect 1491 -138 1493 -136
rect 1495 -138 1497 -136
rect 1469 -145 1471 -143
rect 1473 -145 1475 -143
rect 1469 -146 1475 -145
rect 1482 -144 1486 -142
rect 1482 -146 1483 -144
rect 1485 -146 1486 -144
rect 1491 -143 1497 -138
rect 1491 -145 1493 -143
rect 1495 -145 1497 -143
rect 1491 -146 1497 -145
rect 1523 -138 1525 -136
rect 1527 -138 1529 -136
rect 1523 -143 1529 -138
rect 1545 -138 1547 -136
rect 1549 -138 1551 -136
rect 1523 -145 1525 -143
rect 1527 -145 1529 -143
rect 1523 -146 1529 -145
rect 1534 -144 1538 -142
rect 1534 -146 1535 -144
rect 1537 -146 1538 -144
rect 1545 -143 1551 -138
rect 1580 -138 1582 -136
rect 1584 -138 1586 -136
rect 1580 -139 1586 -138
rect 1621 -138 1623 -136
rect 1625 -138 1627 -136
rect 1621 -139 1627 -138
rect 1545 -145 1547 -143
rect 1549 -145 1551 -143
rect 1545 -146 1551 -145
rect 1602 -143 1619 -142
rect 1602 -145 1604 -143
rect 1606 -145 1619 -143
rect 1602 -146 1619 -145
rect 1650 -143 1656 -136
rect 1650 -145 1652 -143
rect 1654 -145 1656 -143
rect 1650 -146 1656 -145
rect 1661 -143 1665 -141
rect 1661 -145 1662 -143
rect 1664 -145 1665 -143
rect 1403 -148 1409 -147
rect 1394 -152 1395 -150
rect 1397 -151 1398 -150
rect 1397 -152 1411 -151
rect 1394 -155 1411 -152
rect 1345 -176 1363 -175
rect 1345 -178 1347 -176
rect 1349 -178 1363 -176
rect 1345 -179 1363 -178
rect 1407 -167 1411 -155
rect 1407 -169 1408 -167
rect 1410 -169 1411 -167
rect 1407 -174 1411 -169
rect 1399 -178 1411 -174
rect 1399 -182 1403 -178
rect 1414 -181 1415 -179
rect 1285 -185 1286 -183
rect 1288 -184 1310 -183
rect 1288 -185 1306 -184
rect 1285 -186 1306 -185
rect 1308 -186 1310 -184
rect 1176 -187 1201 -186
rect 1285 -187 1310 -186
rect 1315 -187 1319 -185
rect 1383 -183 1403 -182
rect 1383 -185 1385 -183
rect 1387 -185 1403 -183
rect 1383 -186 1403 -185
rect 1439 -150 1463 -146
rect 1482 -150 1486 -146
rect 1437 -154 1443 -150
rect 1459 -151 1499 -150
rect 1459 -153 1483 -151
rect 1485 -153 1499 -151
rect 1437 -164 1441 -154
rect 1447 -155 1451 -153
rect 1459 -154 1499 -153
rect 1447 -157 1448 -155
rect 1450 -157 1451 -155
rect 1447 -158 1451 -157
rect 1437 -166 1438 -164
rect 1440 -166 1441 -164
rect 1437 -168 1441 -166
rect 1444 -162 1451 -158
rect 1444 -173 1448 -162
rect 1487 -167 1491 -162
rect 1487 -169 1488 -167
rect 1490 -169 1491 -167
rect 1430 -174 1448 -173
rect 1430 -176 1432 -174
rect 1434 -175 1448 -174
rect 1434 -176 1459 -175
rect 1430 -177 1455 -176
rect 1444 -178 1455 -177
rect 1457 -178 1459 -176
rect 1444 -179 1459 -178
rect 1464 -176 1468 -174
rect 1464 -178 1465 -176
rect 1467 -178 1468 -176
rect 1464 -183 1468 -178
rect 1487 -171 1491 -169
rect 1495 -165 1499 -154
rect 1495 -167 1501 -165
rect 1495 -169 1498 -167
rect 1500 -169 1501 -167
rect 1495 -171 1501 -169
rect 1495 -174 1499 -171
rect 1479 -178 1499 -174
rect 1479 -182 1483 -178
rect 1443 -184 1465 -183
rect 1434 -187 1438 -185
rect 1443 -186 1445 -184
rect 1447 -185 1465 -184
rect 1467 -185 1468 -183
rect 1447 -186 1468 -185
rect 1473 -183 1483 -182
rect 1473 -185 1475 -183
rect 1477 -185 1483 -183
rect 1473 -186 1483 -185
rect 1534 -150 1538 -146
rect 1557 -150 1581 -146
rect 1521 -151 1561 -150
rect 1521 -153 1535 -151
rect 1537 -153 1561 -151
rect 1521 -154 1561 -153
rect 1521 -165 1525 -154
rect 1569 -155 1573 -153
rect 1577 -154 1583 -150
rect 1569 -157 1570 -155
rect 1572 -157 1573 -155
rect 1569 -158 1573 -157
rect 1569 -162 1576 -158
rect 1519 -167 1525 -165
rect 1519 -169 1520 -167
rect 1522 -169 1525 -167
rect 1519 -171 1525 -169
rect 1529 -167 1533 -162
rect 1529 -169 1530 -167
rect 1532 -169 1533 -167
rect 1529 -171 1533 -169
rect 1521 -174 1525 -171
rect 1521 -178 1541 -174
rect 1537 -182 1541 -178
rect 1572 -173 1576 -162
rect 1579 -164 1583 -154
rect 1579 -166 1580 -164
rect 1582 -166 1583 -164
rect 1579 -168 1583 -166
rect 1572 -174 1590 -173
rect 1552 -176 1556 -174
rect 1572 -175 1586 -174
rect 1552 -178 1553 -176
rect 1555 -178 1556 -176
rect 1537 -183 1547 -182
rect 1537 -185 1543 -183
rect 1545 -185 1547 -183
rect 1537 -186 1547 -185
rect 1552 -183 1556 -178
rect 1561 -176 1586 -175
rect 1588 -176 1590 -174
rect 1561 -178 1563 -176
rect 1565 -177 1590 -176
rect 1565 -178 1576 -177
rect 1561 -179 1576 -178
rect 1615 -150 1619 -146
rect 1615 -154 1630 -150
rect 1605 -163 1611 -162
rect 1626 -167 1630 -154
rect 1633 -157 1634 -146
rect 1626 -169 1627 -167
rect 1629 -169 1630 -167
rect 1626 -175 1630 -169
rect 1661 -150 1665 -145
rect 1670 -145 1676 -136
rect 1701 -138 1703 -136
rect 1705 -138 1707 -136
rect 1701 -139 1707 -138
rect 1736 -138 1738 -136
rect 1740 -138 1742 -136
rect 1670 -147 1672 -145
rect 1674 -147 1676 -145
rect 1736 -143 1742 -138
rect 1758 -138 1760 -136
rect 1762 -138 1764 -136
rect 1736 -145 1738 -143
rect 1740 -145 1742 -143
rect 1736 -146 1742 -145
rect 1749 -144 1753 -142
rect 1749 -146 1750 -144
rect 1752 -146 1753 -144
rect 1758 -143 1764 -138
rect 1758 -145 1760 -143
rect 1762 -145 1764 -143
rect 1758 -146 1764 -145
rect 1790 -138 1792 -136
rect 1794 -138 1796 -136
rect 1790 -143 1796 -138
rect 1812 -138 1814 -136
rect 1816 -138 1818 -136
rect 1790 -145 1792 -143
rect 1794 -145 1796 -143
rect 1790 -146 1796 -145
rect 1801 -144 1805 -142
rect 1801 -146 1802 -144
rect 1804 -146 1805 -144
rect 1812 -143 1818 -138
rect 1847 -138 1849 -136
rect 1851 -138 1853 -136
rect 1847 -139 1853 -138
rect 1888 -138 1890 -136
rect 1892 -138 1894 -136
rect 1888 -139 1894 -138
rect 1931 -138 1932 -136
rect 1934 -138 1935 -136
rect 1812 -145 1814 -143
rect 1816 -145 1818 -143
rect 1812 -146 1818 -145
rect 1869 -143 1886 -142
rect 1869 -145 1871 -143
rect 1873 -145 1886 -143
rect 1869 -146 1886 -145
rect 1670 -148 1676 -147
rect 1661 -152 1662 -150
rect 1664 -151 1665 -150
rect 1664 -152 1678 -151
rect 1661 -155 1678 -152
rect 1612 -176 1630 -175
rect 1612 -178 1614 -176
rect 1616 -178 1630 -176
rect 1612 -179 1630 -178
rect 1674 -167 1678 -155
rect 1674 -169 1675 -167
rect 1677 -169 1678 -167
rect 1674 -174 1678 -169
rect 1666 -178 1678 -174
rect 1666 -182 1670 -178
rect 1681 -181 1682 -179
rect 1552 -185 1553 -183
rect 1555 -184 1577 -183
rect 1555 -185 1573 -184
rect 1552 -186 1573 -185
rect 1575 -186 1577 -184
rect 1443 -187 1468 -186
rect 1552 -187 1577 -186
rect 1582 -187 1586 -185
rect 1650 -183 1670 -182
rect 1650 -185 1652 -183
rect 1654 -185 1670 -183
rect 1650 -186 1670 -185
rect 1706 -150 1730 -146
rect 1749 -150 1753 -146
rect 1704 -154 1710 -150
rect 1726 -151 1766 -150
rect 1726 -153 1750 -151
rect 1752 -153 1766 -151
rect 1704 -164 1708 -154
rect 1714 -155 1718 -153
rect 1726 -154 1766 -153
rect 1714 -157 1715 -155
rect 1717 -157 1718 -155
rect 1714 -158 1718 -157
rect 1704 -166 1705 -164
rect 1707 -166 1708 -164
rect 1704 -168 1708 -166
rect 1711 -162 1718 -158
rect 1711 -173 1715 -162
rect 1754 -167 1758 -162
rect 1754 -169 1755 -167
rect 1757 -169 1758 -167
rect 1697 -174 1715 -173
rect 1697 -176 1699 -174
rect 1701 -175 1715 -174
rect 1701 -176 1726 -175
rect 1697 -177 1722 -176
rect 1711 -178 1722 -177
rect 1724 -178 1726 -176
rect 1711 -179 1726 -178
rect 1731 -176 1735 -174
rect 1731 -178 1732 -176
rect 1734 -178 1735 -176
rect 1731 -183 1735 -178
rect 1754 -171 1758 -169
rect 1762 -165 1766 -154
rect 1762 -167 1768 -165
rect 1762 -169 1765 -167
rect 1767 -169 1768 -167
rect 1762 -171 1768 -169
rect 1762 -174 1766 -171
rect 1746 -178 1766 -174
rect 1746 -182 1750 -178
rect 1710 -184 1732 -183
rect 1701 -187 1705 -185
rect 1710 -186 1712 -184
rect 1714 -185 1732 -184
rect 1734 -185 1735 -183
rect 1714 -186 1735 -185
rect 1740 -183 1750 -182
rect 1740 -185 1742 -183
rect 1744 -185 1750 -183
rect 1740 -186 1750 -185
rect 1801 -150 1805 -146
rect 1824 -150 1848 -146
rect 1788 -151 1828 -150
rect 1788 -153 1802 -151
rect 1804 -153 1828 -151
rect 1788 -154 1828 -153
rect 1788 -165 1792 -154
rect 1836 -155 1840 -153
rect 1844 -154 1850 -150
rect 1836 -157 1837 -155
rect 1839 -157 1840 -155
rect 1836 -158 1840 -157
rect 1836 -162 1843 -158
rect 1786 -167 1792 -165
rect 1786 -169 1787 -167
rect 1789 -169 1792 -167
rect 1786 -171 1792 -169
rect 1796 -167 1800 -162
rect 1796 -169 1797 -167
rect 1799 -169 1800 -167
rect 1796 -171 1800 -169
rect 1788 -174 1792 -171
rect 1788 -178 1808 -174
rect 1804 -182 1808 -178
rect 1839 -173 1843 -162
rect 1846 -164 1850 -154
rect 1846 -166 1847 -164
rect 1849 -166 1850 -164
rect 1846 -168 1850 -166
rect 1839 -174 1857 -173
rect 1819 -176 1823 -174
rect 1839 -175 1853 -174
rect 1819 -178 1820 -176
rect 1822 -178 1823 -176
rect 1804 -183 1814 -182
rect 1804 -185 1810 -183
rect 1812 -185 1814 -183
rect 1804 -186 1814 -185
rect 1819 -183 1823 -178
rect 1828 -176 1853 -175
rect 1855 -176 1857 -174
rect 1828 -178 1830 -176
rect 1832 -177 1857 -176
rect 1882 -150 1886 -146
rect 1882 -154 1897 -150
rect 1872 -163 1878 -162
rect 1893 -167 1897 -154
rect 1900 -157 1901 -146
rect 1893 -169 1894 -167
rect 1896 -169 1897 -167
rect 1893 -175 1897 -169
rect 1931 -143 1935 -138
rect 1987 -138 1989 -136
rect 1991 -138 1993 -136
rect 1987 -139 1993 -138
rect 2022 -138 2024 -136
rect 2026 -138 2028 -136
rect 1931 -145 1932 -143
rect 1934 -145 1935 -143
rect 1931 -147 1935 -145
rect 1939 -142 1972 -141
rect 1939 -144 1968 -142
rect 1970 -144 1972 -142
rect 1939 -145 1972 -144
rect 2022 -143 2028 -138
rect 2044 -138 2046 -136
rect 2048 -138 2050 -136
rect 2022 -145 2024 -143
rect 2026 -145 2028 -143
rect 1939 -156 1943 -145
rect 2022 -146 2028 -145
rect 2035 -144 2039 -142
rect 2035 -146 2036 -144
rect 2038 -146 2039 -144
rect 2044 -143 2050 -138
rect 2044 -145 2046 -143
rect 2048 -145 2050 -143
rect 2044 -146 2050 -145
rect 2076 -138 2078 -136
rect 2080 -138 2082 -136
rect 2076 -143 2082 -138
rect 2098 -138 2100 -136
rect 2102 -138 2104 -136
rect 2076 -145 2078 -143
rect 2080 -145 2082 -143
rect 2076 -146 2082 -145
rect 2087 -144 2091 -142
rect 2087 -146 2088 -144
rect 2090 -146 2091 -144
rect 2098 -143 2104 -138
rect 2133 -138 2135 -136
rect 2137 -138 2139 -136
rect 2133 -139 2139 -138
rect 2174 -138 2176 -136
rect 2178 -138 2180 -136
rect 2174 -139 2180 -138
rect 2210 -138 2211 -136
rect 2213 -138 2214 -136
rect 2210 -140 2214 -138
rect 2243 -138 2245 -136
rect 2247 -138 2249 -136
rect 2243 -139 2249 -138
rect 2278 -138 2279 -136
rect 2281 -138 2282 -136
rect 2278 -140 2282 -138
rect 2311 -138 2313 -136
rect 2315 -138 2317 -136
rect 2311 -139 2317 -138
rect 2098 -145 2100 -143
rect 2102 -145 2104 -143
rect 2098 -146 2104 -145
rect 2155 -143 2172 -142
rect 2155 -145 2157 -143
rect 2159 -145 2172 -143
rect 2155 -146 2172 -145
rect 1920 -157 1943 -156
rect 1920 -159 1922 -157
rect 1924 -159 1943 -157
rect 1920 -160 1943 -159
rect 1920 -166 1924 -160
rect 1832 -178 1843 -177
rect 1828 -179 1843 -178
rect 1879 -176 1897 -175
rect 1879 -178 1881 -176
rect 1883 -178 1897 -176
rect 1879 -179 1897 -178
rect 1913 -170 1924 -166
rect 1913 -176 1917 -170
rect 1939 -166 1943 -160
rect 1947 -150 1951 -148
rect 1947 -152 1948 -150
rect 1950 -152 1951 -150
rect 1947 -157 1951 -152
rect 1947 -159 1948 -157
rect 1950 -158 1951 -157
rect 1950 -159 1963 -158
rect 1947 -162 1963 -159
rect 1959 -164 1963 -162
rect 1959 -166 1964 -164
rect 1939 -167 1955 -166
rect 1939 -169 1951 -167
rect 1953 -169 1955 -167
rect 1939 -170 1955 -169
rect 1959 -168 1961 -166
rect 1963 -168 1964 -166
rect 1959 -170 1964 -168
rect 1913 -178 1914 -176
rect 1916 -178 1917 -176
rect 1913 -180 1917 -178
rect 1959 -174 1963 -170
rect 1939 -178 1963 -174
rect 1939 -181 1943 -178
rect 1939 -183 1940 -181
rect 1942 -183 1943 -181
rect 1819 -185 1820 -183
rect 1822 -184 1844 -183
rect 1822 -185 1840 -184
rect 1819 -186 1840 -185
rect 1842 -186 1844 -184
rect 1710 -187 1735 -186
rect 1819 -187 1844 -186
rect 1849 -187 1853 -185
rect 1926 -184 1932 -183
rect 1926 -186 1928 -184
rect 1930 -186 1932 -184
rect 1939 -185 1943 -183
rect 1992 -150 2016 -146
rect 2035 -150 2039 -146
rect 1990 -154 1996 -150
rect 2012 -151 2052 -150
rect 2012 -153 2036 -151
rect 2038 -153 2052 -151
rect 1990 -164 1994 -154
rect 2000 -155 2004 -153
rect 2012 -154 2052 -153
rect 2000 -157 2001 -155
rect 2003 -157 2004 -155
rect 2000 -158 2004 -157
rect 1990 -166 1991 -164
rect 1993 -166 1994 -164
rect 1990 -168 1994 -166
rect 1997 -162 2004 -158
rect 1997 -173 2001 -162
rect 2040 -167 2044 -162
rect 2040 -169 2041 -167
rect 2043 -169 2044 -167
rect 1983 -174 2001 -173
rect 1983 -176 1985 -174
rect 1987 -175 2001 -174
rect 1987 -176 2012 -175
rect 1983 -177 2008 -176
rect 1997 -178 2008 -177
rect 2010 -178 2012 -176
rect 1997 -179 2012 -178
rect 2017 -176 2021 -174
rect 2017 -178 2018 -176
rect 2020 -178 2021 -176
rect 2017 -183 2021 -178
rect 2040 -171 2044 -169
rect 2048 -165 2052 -154
rect 2048 -167 2054 -165
rect 2048 -169 2051 -167
rect 2053 -169 2054 -167
rect 2048 -171 2054 -169
rect 2048 -174 2052 -171
rect 2032 -178 2052 -174
rect 2032 -182 2036 -178
rect 1996 -184 2018 -183
rect 99 -189 100 -187
rect 102 -189 103 -187
rect 247 -189 248 -187
rect 250 -189 251 -187
rect 99 -192 103 -189
rect 155 -190 161 -189
rect 155 -192 157 -190
rect 159 -192 161 -190
rect 189 -190 195 -189
rect 189 -192 191 -190
rect 193 -192 195 -190
rect 247 -192 251 -189
rect 267 -189 273 -188
rect 267 -191 269 -189
rect 271 -191 273 -189
rect 267 -192 273 -191
rect 286 -189 292 -188
rect 286 -191 288 -189
rect 290 -191 292 -189
rect 286 -192 292 -191
rect 366 -189 367 -187
rect 369 -189 370 -187
rect 514 -189 515 -187
rect 517 -189 518 -187
rect 366 -192 370 -189
rect 422 -190 428 -189
rect 422 -192 424 -190
rect 426 -192 428 -190
rect 456 -190 462 -189
rect 456 -192 458 -190
rect 460 -192 462 -190
rect 514 -192 518 -189
rect 534 -189 540 -188
rect 534 -191 536 -189
rect 538 -191 540 -189
rect 534 -192 540 -191
rect 553 -189 559 -188
rect 553 -191 555 -189
rect 557 -191 559 -189
rect 553 -192 559 -191
rect 633 -189 634 -187
rect 636 -189 637 -187
rect 781 -189 782 -187
rect 784 -189 785 -187
rect 633 -192 637 -189
rect 689 -190 695 -189
rect 689 -192 691 -190
rect 693 -192 695 -190
rect 723 -190 729 -189
rect 723 -192 725 -190
rect 727 -192 729 -190
rect 781 -192 785 -189
rect 801 -189 807 -188
rect 801 -191 803 -189
rect 805 -191 807 -189
rect 801 -192 807 -191
rect 820 -189 826 -188
rect 820 -191 822 -189
rect 824 -191 826 -189
rect 820 -192 826 -191
rect 900 -189 901 -187
rect 903 -189 904 -187
rect 1048 -189 1049 -187
rect 1051 -189 1052 -187
rect 900 -192 904 -189
rect 956 -190 962 -189
rect 956 -192 958 -190
rect 960 -192 962 -190
rect 990 -190 996 -189
rect 990 -192 992 -190
rect 994 -192 996 -190
rect 1048 -192 1052 -189
rect 1068 -189 1074 -188
rect 1068 -191 1070 -189
rect 1072 -191 1074 -189
rect 1068 -192 1074 -191
rect 1087 -189 1093 -188
rect 1087 -191 1089 -189
rect 1091 -191 1093 -189
rect 1087 -192 1093 -191
rect 1167 -189 1168 -187
rect 1170 -189 1171 -187
rect 1315 -189 1316 -187
rect 1318 -189 1319 -187
rect 1167 -192 1171 -189
rect 1223 -190 1229 -189
rect 1223 -192 1225 -190
rect 1227 -192 1229 -190
rect 1257 -190 1263 -189
rect 1257 -192 1259 -190
rect 1261 -192 1263 -190
rect 1315 -192 1319 -189
rect 1335 -189 1341 -188
rect 1335 -191 1337 -189
rect 1339 -191 1341 -189
rect 1335 -192 1341 -191
rect 1354 -189 1360 -188
rect 1354 -191 1356 -189
rect 1358 -191 1360 -189
rect 1354 -192 1360 -191
rect 1434 -189 1435 -187
rect 1437 -189 1438 -187
rect 1582 -189 1583 -187
rect 1585 -189 1586 -187
rect 1434 -192 1438 -189
rect 1490 -190 1496 -189
rect 1490 -192 1492 -190
rect 1494 -192 1496 -190
rect 1524 -190 1530 -189
rect 1524 -192 1526 -190
rect 1528 -192 1530 -190
rect 1582 -192 1586 -189
rect 1602 -189 1608 -188
rect 1602 -191 1604 -189
rect 1606 -191 1608 -189
rect 1602 -192 1608 -191
rect 1621 -189 1627 -188
rect 1621 -191 1623 -189
rect 1625 -191 1627 -189
rect 1621 -192 1627 -191
rect 1701 -189 1702 -187
rect 1704 -189 1705 -187
rect 1849 -189 1850 -187
rect 1852 -189 1853 -187
rect 1701 -192 1705 -189
rect 1757 -190 1763 -189
rect 1757 -192 1759 -190
rect 1761 -192 1763 -190
rect 1791 -190 1797 -189
rect 1791 -192 1793 -190
rect 1795 -192 1797 -190
rect 1849 -192 1853 -189
rect 1869 -189 1875 -188
rect 1869 -191 1871 -189
rect 1873 -191 1875 -189
rect 1869 -192 1875 -191
rect 1888 -189 1894 -188
rect 1888 -191 1890 -189
rect 1892 -191 1894 -189
rect 1888 -192 1894 -191
rect 1926 -192 1932 -186
rect 1987 -187 1991 -185
rect 1996 -186 1998 -184
rect 2000 -185 2018 -184
rect 2020 -185 2021 -183
rect 2000 -186 2021 -185
rect 2026 -183 2036 -182
rect 2026 -185 2028 -183
rect 2030 -185 2036 -183
rect 2026 -186 2036 -185
rect 2087 -150 2091 -146
rect 2110 -150 2134 -146
rect 2074 -151 2114 -150
rect 2074 -153 2088 -151
rect 2090 -153 2114 -151
rect 2074 -154 2114 -153
rect 2074 -165 2078 -154
rect 2122 -155 2126 -153
rect 2130 -154 2136 -150
rect 2122 -157 2123 -155
rect 2125 -157 2126 -155
rect 2122 -158 2126 -157
rect 2122 -162 2129 -158
rect 2072 -167 2078 -165
rect 2072 -169 2073 -167
rect 2075 -169 2078 -167
rect 2072 -171 2078 -169
rect 2082 -167 2086 -162
rect 2082 -169 2083 -167
rect 2085 -169 2086 -167
rect 2082 -171 2086 -169
rect 2074 -174 2078 -171
rect 2074 -178 2094 -174
rect 2090 -182 2094 -178
rect 2125 -173 2129 -162
rect 2132 -164 2136 -154
rect 2132 -166 2133 -164
rect 2135 -166 2136 -164
rect 2132 -168 2136 -166
rect 2125 -174 2143 -173
rect 2105 -176 2109 -174
rect 2125 -175 2139 -174
rect 2105 -178 2106 -176
rect 2108 -178 2109 -176
rect 2090 -183 2100 -182
rect 2090 -185 2096 -183
rect 2098 -185 2100 -183
rect 2090 -186 2100 -185
rect 2105 -183 2109 -178
rect 2114 -176 2139 -175
rect 2141 -176 2143 -174
rect 2114 -178 2116 -176
rect 2118 -177 2143 -176
rect 2118 -178 2129 -177
rect 2114 -179 2129 -178
rect 2168 -150 2172 -146
rect 2168 -154 2183 -150
rect 2158 -163 2164 -162
rect 2179 -167 2183 -154
rect 2186 -157 2187 -146
rect 2226 -146 2239 -145
rect 2226 -148 2228 -146
rect 2230 -148 2239 -146
rect 2226 -149 2239 -148
rect 2235 -153 2251 -149
rect 2179 -169 2180 -167
rect 2182 -169 2183 -167
rect 2179 -175 2183 -169
rect 2223 -157 2227 -155
rect 2165 -176 2183 -175
rect 2165 -178 2167 -176
rect 2169 -178 2183 -176
rect 2165 -179 2183 -178
rect 2199 -158 2224 -157
rect 2199 -160 2201 -158
rect 2203 -159 2224 -158
rect 2226 -159 2227 -157
rect 2203 -160 2227 -159
rect 2199 -161 2227 -160
rect 2105 -185 2106 -183
rect 2108 -184 2130 -183
rect 2108 -185 2126 -184
rect 2105 -186 2126 -185
rect 2128 -186 2130 -184
rect 2199 -181 2203 -161
rect 2223 -171 2227 -161
rect 2243 -166 2244 -160
rect 2247 -170 2251 -153
rect 2223 -173 2234 -171
rect 2223 -175 2231 -173
rect 2233 -175 2234 -173
rect 2247 -172 2252 -170
rect 2247 -174 2249 -172
rect 2251 -174 2252 -172
rect 2223 -177 2234 -175
rect 2237 -176 2252 -174
rect 2237 -178 2251 -176
rect 2199 -182 2205 -181
rect 2199 -184 2201 -182
rect 2203 -184 2205 -182
rect 2199 -185 2205 -184
rect 2209 -182 2215 -181
rect 2209 -184 2211 -182
rect 2213 -184 2215 -182
rect 2237 -183 2241 -178
rect 2294 -146 2307 -145
rect 2294 -148 2296 -146
rect 2298 -148 2307 -146
rect 2294 -149 2307 -148
rect 2303 -153 2319 -149
rect 2291 -157 2295 -155
rect 1996 -187 2021 -186
rect 2105 -187 2130 -186
rect 2135 -187 2139 -185
rect 1987 -189 1988 -187
rect 1990 -189 1991 -187
rect 2135 -189 2136 -187
rect 2138 -189 2139 -187
rect 1987 -192 1991 -189
rect 2043 -190 2049 -189
rect 2043 -192 2045 -190
rect 2047 -192 2049 -190
rect 2077 -190 2083 -189
rect 2077 -192 2079 -190
rect 2081 -192 2083 -190
rect 2135 -192 2139 -189
rect 2155 -189 2161 -188
rect 2155 -191 2157 -189
rect 2159 -191 2161 -189
rect 2155 -192 2161 -191
rect 2174 -189 2180 -188
rect 2174 -191 2176 -189
rect 2178 -191 2180 -189
rect 2174 -192 2180 -191
rect 2209 -192 2215 -184
rect 2226 -184 2241 -183
rect 2226 -186 2228 -184
rect 2230 -186 2241 -184
rect 2226 -187 2241 -186
rect 2244 -184 2248 -182
rect 2244 -186 2245 -184
rect 2247 -186 2248 -184
rect 2267 -158 2292 -157
rect 2267 -160 2269 -158
rect 2271 -159 2292 -158
rect 2294 -159 2295 -157
rect 2271 -160 2295 -159
rect 2267 -161 2295 -160
rect 2267 -181 2271 -161
rect 2291 -171 2295 -161
rect 2311 -166 2312 -160
rect 2315 -170 2319 -153
rect 2291 -173 2302 -171
rect 2291 -175 2299 -173
rect 2301 -175 2302 -173
rect 2315 -172 2320 -170
rect 2315 -174 2317 -172
rect 2319 -174 2320 -172
rect 2291 -177 2302 -175
rect 2305 -176 2320 -174
rect 2305 -178 2319 -176
rect 2267 -182 2273 -181
rect 2267 -184 2269 -182
rect 2271 -184 2273 -182
rect 2267 -185 2273 -184
rect 2277 -182 2283 -181
rect 2277 -184 2279 -182
rect 2281 -184 2283 -182
rect 2305 -183 2309 -178
rect 2244 -192 2248 -186
rect 2277 -192 2283 -184
rect 2294 -184 2309 -183
rect 2294 -186 2296 -184
rect 2298 -186 2309 -184
rect 2294 -187 2309 -186
rect 2312 -184 2316 -182
rect 2312 -186 2313 -184
rect 2315 -186 2316 -184
rect 2312 -192 2316 -186
rect 99 -211 103 -208
rect 155 -210 157 -208
rect 159 -210 161 -208
rect 155 -211 161 -210
rect 189 -210 191 -208
rect 193 -210 195 -208
rect 189 -211 195 -210
rect 247 -211 251 -208
rect 99 -213 100 -211
rect 102 -213 103 -211
rect 247 -213 248 -211
rect 250 -213 251 -211
rect 267 -209 273 -208
rect 267 -211 269 -209
rect 271 -211 273 -209
rect 267 -212 273 -211
rect 286 -209 292 -208
rect 286 -211 288 -209
rect 290 -211 292 -209
rect 286 -212 292 -211
rect 366 -211 370 -208
rect 422 -210 424 -208
rect 426 -210 428 -208
rect 422 -211 428 -210
rect 456 -210 458 -208
rect 460 -210 462 -208
rect 456 -211 462 -210
rect 514 -211 518 -208
rect 366 -213 367 -211
rect 369 -213 370 -211
rect 514 -213 515 -211
rect 517 -213 518 -211
rect 534 -209 540 -208
rect 534 -211 536 -209
rect 538 -211 540 -209
rect 534 -212 540 -211
rect 553 -209 559 -208
rect 553 -211 555 -209
rect 557 -211 559 -209
rect 553 -212 559 -211
rect 633 -211 637 -208
rect 689 -210 691 -208
rect 693 -210 695 -208
rect 689 -211 695 -210
rect 723 -210 725 -208
rect 727 -210 729 -208
rect 723 -211 729 -210
rect 781 -211 785 -208
rect 633 -213 634 -211
rect 636 -213 637 -211
rect 781 -213 782 -211
rect 784 -213 785 -211
rect 801 -209 807 -208
rect 801 -211 803 -209
rect 805 -211 807 -209
rect 801 -212 807 -211
rect 820 -209 826 -208
rect 820 -211 822 -209
rect 824 -211 826 -209
rect 820 -212 826 -211
rect 900 -211 904 -208
rect 956 -210 958 -208
rect 960 -210 962 -208
rect 956 -211 962 -210
rect 990 -210 992 -208
rect 994 -210 996 -208
rect 990 -211 996 -210
rect 1048 -211 1052 -208
rect 900 -213 901 -211
rect 903 -213 904 -211
rect 1048 -213 1049 -211
rect 1051 -213 1052 -211
rect 1068 -209 1074 -208
rect 1068 -211 1070 -209
rect 1072 -211 1074 -209
rect 1068 -212 1074 -211
rect 1087 -209 1093 -208
rect 1087 -211 1089 -209
rect 1091 -211 1093 -209
rect 1087 -212 1093 -211
rect 1167 -211 1171 -208
rect 1223 -210 1225 -208
rect 1227 -210 1229 -208
rect 1223 -211 1229 -210
rect 1257 -210 1259 -208
rect 1261 -210 1263 -208
rect 1257 -211 1263 -210
rect 1315 -211 1319 -208
rect 1167 -213 1168 -211
rect 1170 -213 1171 -211
rect 1315 -213 1316 -211
rect 1318 -213 1319 -211
rect 1335 -209 1341 -208
rect 1335 -211 1337 -209
rect 1339 -211 1341 -209
rect 1335 -212 1341 -211
rect 1354 -209 1360 -208
rect 1354 -211 1356 -209
rect 1358 -211 1360 -209
rect 1354 -212 1360 -211
rect 1434 -211 1438 -208
rect 1490 -210 1492 -208
rect 1494 -210 1496 -208
rect 1490 -211 1496 -210
rect 1524 -210 1526 -208
rect 1528 -210 1530 -208
rect 1524 -211 1530 -210
rect 1582 -211 1586 -208
rect 1434 -213 1435 -211
rect 1437 -213 1438 -211
rect 1582 -213 1583 -211
rect 1585 -213 1586 -211
rect 1602 -209 1608 -208
rect 1602 -211 1604 -209
rect 1606 -211 1608 -209
rect 1602 -212 1608 -211
rect 1621 -209 1627 -208
rect 1621 -211 1623 -209
rect 1625 -211 1627 -209
rect 1621 -212 1627 -211
rect 1701 -211 1705 -208
rect 1757 -210 1759 -208
rect 1761 -210 1763 -208
rect 1757 -211 1763 -210
rect 1791 -210 1793 -208
rect 1795 -210 1797 -208
rect 1791 -211 1797 -210
rect 1849 -211 1853 -208
rect 1701 -213 1702 -211
rect 1704 -213 1705 -211
rect 1849 -213 1850 -211
rect 1852 -213 1853 -211
rect 1869 -209 1875 -208
rect 1869 -211 1871 -209
rect 1873 -211 1875 -209
rect 1869 -212 1875 -211
rect 1888 -209 1894 -208
rect 1888 -211 1890 -209
rect 1892 -211 1894 -209
rect 1888 -212 1894 -211
rect 8 -215 28 -214
rect 8 -217 10 -215
rect 12 -217 28 -215
rect 8 -218 28 -217
rect 24 -222 28 -218
rect 48 -215 68 -214
rect 48 -217 50 -215
rect 52 -217 68 -215
rect 48 -218 68 -217
rect 39 -221 40 -219
rect 24 -226 36 -222
rect 32 -231 36 -226
rect 32 -233 33 -231
rect 35 -233 36 -231
rect 32 -245 36 -233
rect 64 -222 68 -218
rect 79 -221 80 -219
rect 64 -226 76 -222
rect 72 -231 76 -226
rect 72 -233 73 -231
rect 75 -233 76 -231
rect 19 -248 36 -245
rect 19 -250 20 -248
rect 22 -249 36 -248
rect 22 -250 23 -249
rect 8 -255 14 -254
rect 8 -257 10 -255
rect 12 -257 14 -255
rect 8 -264 14 -257
rect 19 -255 23 -250
rect 72 -245 76 -233
rect 59 -248 76 -245
rect 59 -250 60 -248
rect 62 -249 76 -248
rect 62 -250 63 -249
rect 19 -257 20 -255
rect 22 -257 23 -255
rect 19 -259 23 -257
rect 28 -253 34 -252
rect 28 -255 30 -253
rect 32 -255 34 -253
rect 28 -264 34 -255
rect 48 -255 54 -254
rect 48 -257 50 -255
rect 52 -257 54 -255
rect 48 -264 54 -257
rect 59 -255 63 -250
rect 99 -215 103 -213
rect 108 -214 133 -213
rect 217 -214 242 -213
rect 108 -216 110 -214
rect 112 -215 133 -214
rect 112 -216 130 -215
rect 108 -217 130 -216
rect 132 -217 133 -215
rect 109 -222 124 -221
rect 109 -223 120 -222
rect 95 -224 120 -223
rect 122 -224 124 -222
rect 95 -226 97 -224
rect 99 -225 124 -224
rect 129 -222 133 -217
rect 138 -215 148 -214
rect 138 -217 140 -215
rect 142 -217 148 -215
rect 138 -218 148 -217
rect 129 -224 130 -222
rect 132 -224 133 -222
rect 99 -226 113 -225
rect 129 -226 133 -224
rect 95 -227 113 -226
rect 102 -234 106 -232
rect 102 -236 103 -234
rect 105 -236 106 -234
rect 102 -246 106 -236
rect 109 -238 113 -227
rect 144 -222 148 -218
rect 144 -226 164 -222
rect 160 -229 164 -226
rect 152 -231 156 -229
rect 152 -233 153 -231
rect 155 -233 156 -231
rect 152 -238 156 -233
rect 160 -231 166 -229
rect 160 -233 163 -231
rect 165 -233 166 -231
rect 160 -235 166 -233
rect 109 -242 116 -238
rect 112 -243 116 -242
rect 112 -245 113 -243
rect 115 -245 116 -243
rect 102 -250 108 -246
rect 112 -247 116 -245
rect 160 -246 164 -235
rect 124 -247 164 -246
rect 124 -249 148 -247
rect 150 -249 164 -247
rect 124 -250 164 -249
rect 59 -257 60 -255
rect 62 -257 63 -255
rect 59 -259 63 -257
rect 68 -253 74 -252
rect 68 -255 70 -253
rect 72 -255 74 -253
rect 104 -254 128 -250
rect 147 -254 151 -250
rect 202 -215 212 -214
rect 202 -217 208 -215
rect 210 -217 212 -215
rect 202 -218 212 -217
rect 217 -215 238 -214
rect 217 -217 218 -215
rect 220 -216 238 -215
rect 240 -216 242 -214
rect 247 -215 251 -213
rect 220 -217 242 -216
rect 202 -222 206 -218
rect 186 -226 206 -222
rect 186 -229 190 -226
rect 184 -231 190 -229
rect 184 -233 185 -231
rect 187 -233 190 -231
rect 184 -235 190 -233
rect 186 -246 190 -235
rect 194 -231 198 -229
rect 217 -222 221 -217
rect 315 -215 335 -214
rect 315 -217 317 -215
rect 319 -217 335 -215
rect 315 -218 335 -217
rect 217 -224 218 -222
rect 220 -224 221 -222
rect 217 -226 221 -224
rect 226 -222 241 -221
rect 226 -224 228 -222
rect 230 -223 241 -222
rect 230 -224 255 -223
rect 226 -225 251 -224
rect 237 -226 251 -225
rect 253 -226 255 -224
rect 237 -227 255 -226
rect 194 -233 195 -231
rect 197 -233 198 -231
rect 194 -238 198 -233
rect 237 -238 241 -227
rect 234 -242 241 -238
rect 244 -234 248 -232
rect 244 -236 245 -234
rect 247 -236 248 -234
rect 234 -243 238 -242
rect 234 -245 235 -243
rect 237 -245 238 -243
rect 186 -247 226 -246
rect 234 -247 238 -245
rect 244 -246 248 -236
rect 277 -222 295 -221
rect 277 -224 279 -222
rect 281 -224 295 -222
rect 277 -225 295 -224
rect 291 -231 295 -225
rect 291 -233 292 -231
rect 294 -233 295 -231
rect 270 -238 276 -237
rect 186 -249 200 -247
rect 202 -249 226 -247
rect 186 -250 226 -249
rect 242 -250 248 -246
rect 199 -254 203 -250
rect 222 -254 246 -250
rect 291 -246 295 -233
rect 280 -250 295 -246
rect 280 -254 284 -250
rect 298 -254 299 -243
rect 331 -222 335 -218
rect 346 -221 347 -219
rect 331 -226 343 -222
rect 339 -231 343 -226
rect 339 -233 340 -231
rect 342 -233 343 -231
rect 339 -245 343 -233
rect 326 -248 343 -245
rect 326 -250 327 -248
rect 329 -249 343 -248
rect 329 -250 330 -249
rect 68 -264 74 -255
rect 134 -255 140 -254
rect 134 -257 136 -255
rect 138 -257 140 -255
rect 99 -262 105 -261
rect 99 -264 101 -262
rect 103 -264 105 -262
rect 134 -262 140 -257
rect 147 -256 148 -254
rect 150 -256 151 -254
rect 147 -258 151 -256
rect 156 -255 162 -254
rect 156 -257 158 -255
rect 160 -257 162 -255
rect 134 -264 136 -262
rect 138 -264 140 -262
rect 156 -262 162 -257
rect 156 -264 158 -262
rect 160 -264 162 -262
rect 188 -255 194 -254
rect 188 -257 190 -255
rect 192 -257 194 -255
rect 188 -262 194 -257
rect 199 -256 200 -254
rect 202 -256 203 -254
rect 199 -258 203 -256
rect 210 -255 216 -254
rect 210 -257 212 -255
rect 214 -257 216 -255
rect 188 -264 190 -262
rect 192 -264 194 -262
rect 210 -262 216 -257
rect 267 -255 284 -254
rect 267 -257 269 -255
rect 271 -257 284 -255
rect 267 -258 284 -257
rect 315 -255 321 -254
rect 315 -257 317 -255
rect 319 -257 321 -255
rect 210 -264 212 -262
rect 214 -264 216 -262
rect 245 -262 251 -261
rect 245 -264 247 -262
rect 249 -264 251 -262
rect 286 -262 292 -261
rect 286 -264 288 -262
rect 290 -264 292 -262
rect 315 -264 321 -257
rect 326 -255 330 -250
rect 366 -215 370 -213
rect 375 -214 400 -213
rect 484 -214 509 -213
rect 375 -216 377 -214
rect 379 -215 400 -214
rect 379 -216 397 -215
rect 375 -217 397 -216
rect 399 -217 400 -215
rect 376 -222 391 -221
rect 376 -223 387 -222
rect 362 -224 387 -223
rect 389 -224 391 -222
rect 362 -226 364 -224
rect 366 -225 391 -224
rect 396 -222 400 -217
rect 405 -215 415 -214
rect 405 -217 407 -215
rect 409 -217 415 -215
rect 405 -218 415 -217
rect 396 -224 397 -222
rect 399 -224 400 -222
rect 366 -226 380 -225
rect 396 -226 400 -224
rect 362 -227 380 -226
rect 369 -234 373 -232
rect 369 -236 370 -234
rect 372 -236 373 -234
rect 369 -246 373 -236
rect 376 -238 380 -227
rect 411 -222 415 -218
rect 411 -226 431 -222
rect 427 -229 431 -226
rect 419 -231 423 -229
rect 419 -233 420 -231
rect 422 -233 423 -231
rect 419 -238 423 -233
rect 427 -231 433 -229
rect 427 -233 430 -231
rect 432 -233 433 -231
rect 427 -235 433 -233
rect 376 -242 383 -238
rect 379 -243 383 -242
rect 379 -245 380 -243
rect 382 -245 383 -243
rect 369 -250 375 -246
rect 379 -247 383 -245
rect 427 -246 431 -235
rect 391 -247 431 -246
rect 391 -249 415 -247
rect 417 -249 431 -247
rect 391 -250 431 -249
rect 326 -257 327 -255
rect 329 -257 330 -255
rect 326 -259 330 -257
rect 335 -253 341 -252
rect 335 -255 337 -253
rect 339 -255 341 -253
rect 371 -254 395 -250
rect 414 -254 418 -250
rect 469 -215 479 -214
rect 469 -217 475 -215
rect 477 -217 479 -215
rect 469 -218 479 -217
rect 484 -215 505 -214
rect 484 -217 485 -215
rect 487 -216 505 -215
rect 507 -216 509 -214
rect 514 -215 518 -213
rect 487 -217 509 -216
rect 469 -222 473 -218
rect 453 -226 473 -222
rect 453 -229 457 -226
rect 451 -231 457 -229
rect 451 -233 452 -231
rect 454 -233 457 -231
rect 451 -235 457 -233
rect 453 -246 457 -235
rect 461 -231 465 -229
rect 484 -222 488 -217
rect 582 -215 602 -214
rect 582 -217 584 -215
rect 586 -217 602 -215
rect 582 -218 602 -217
rect 484 -224 485 -222
rect 487 -224 488 -222
rect 484 -226 488 -224
rect 493 -222 508 -221
rect 493 -224 495 -222
rect 497 -223 508 -222
rect 497 -224 522 -223
rect 493 -225 518 -224
rect 504 -226 518 -225
rect 520 -226 522 -224
rect 504 -227 522 -226
rect 461 -233 462 -231
rect 464 -233 465 -231
rect 461 -238 465 -233
rect 504 -238 508 -227
rect 501 -242 508 -238
rect 511 -234 515 -232
rect 511 -236 512 -234
rect 514 -236 515 -234
rect 501 -243 505 -242
rect 501 -245 502 -243
rect 504 -245 505 -243
rect 453 -247 493 -246
rect 501 -247 505 -245
rect 511 -246 515 -236
rect 544 -222 562 -221
rect 544 -224 546 -222
rect 548 -224 562 -222
rect 544 -225 562 -224
rect 558 -231 562 -225
rect 558 -233 559 -231
rect 561 -233 562 -231
rect 537 -238 543 -237
rect 453 -249 467 -247
rect 469 -249 493 -247
rect 453 -250 493 -249
rect 509 -250 515 -246
rect 466 -254 470 -250
rect 489 -254 513 -250
rect 558 -246 562 -233
rect 547 -250 562 -246
rect 547 -254 551 -250
rect 565 -254 566 -243
rect 598 -222 602 -218
rect 613 -221 614 -219
rect 598 -226 610 -222
rect 606 -231 610 -226
rect 606 -233 607 -231
rect 609 -233 610 -231
rect 606 -245 610 -233
rect 593 -248 610 -245
rect 593 -250 594 -248
rect 596 -249 610 -248
rect 596 -250 597 -249
rect 335 -264 341 -255
rect 401 -255 407 -254
rect 401 -257 403 -255
rect 405 -257 407 -255
rect 366 -262 372 -261
rect 366 -264 368 -262
rect 370 -264 372 -262
rect 401 -262 407 -257
rect 414 -256 415 -254
rect 417 -256 418 -254
rect 414 -258 418 -256
rect 423 -255 429 -254
rect 423 -257 425 -255
rect 427 -257 429 -255
rect 401 -264 403 -262
rect 405 -264 407 -262
rect 423 -262 429 -257
rect 423 -264 425 -262
rect 427 -264 429 -262
rect 455 -255 461 -254
rect 455 -257 457 -255
rect 459 -257 461 -255
rect 455 -262 461 -257
rect 466 -256 467 -254
rect 469 -256 470 -254
rect 466 -258 470 -256
rect 477 -255 483 -254
rect 477 -257 479 -255
rect 481 -257 483 -255
rect 455 -264 457 -262
rect 459 -264 461 -262
rect 477 -262 483 -257
rect 534 -255 551 -254
rect 534 -257 536 -255
rect 538 -257 551 -255
rect 534 -258 551 -257
rect 582 -255 588 -254
rect 582 -257 584 -255
rect 586 -257 588 -255
rect 477 -264 479 -262
rect 481 -264 483 -262
rect 512 -262 518 -261
rect 512 -264 514 -262
rect 516 -264 518 -262
rect 553 -262 559 -261
rect 553 -264 555 -262
rect 557 -264 559 -262
rect 582 -264 588 -257
rect 593 -255 597 -250
rect 633 -215 637 -213
rect 642 -214 667 -213
rect 751 -214 776 -213
rect 642 -216 644 -214
rect 646 -215 667 -214
rect 646 -216 664 -215
rect 642 -217 664 -216
rect 666 -217 667 -215
rect 643 -222 658 -221
rect 643 -223 654 -222
rect 629 -224 654 -223
rect 656 -224 658 -222
rect 629 -226 631 -224
rect 633 -225 658 -224
rect 663 -222 667 -217
rect 672 -215 682 -214
rect 672 -217 674 -215
rect 676 -217 682 -215
rect 672 -218 682 -217
rect 663 -224 664 -222
rect 666 -224 667 -222
rect 633 -226 647 -225
rect 663 -226 667 -224
rect 629 -227 647 -226
rect 636 -234 640 -232
rect 636 -236 637 -234
rect 639 -236 640 -234
rect 636 -246 640 -236
rect 643 -238 647 -227
rect 678 -222 682 -218
rect 678 -226 698 -222
rect 694 -229 698 -226
rect 686 -231 690 -229
rect 686 -233 687 -231
rect 689 -233 690 -231
rect 686 -238 690 -233
rect 694 -231 700 -229
rect 694 -233 697 -231
rect 699 -233 700 -231
rect 694 -235 700 -233
rect 643 -242 650 -238
rect 646 -243 650 -242
rect 646 -245 647 -243
rect 649 -245 650 -243
rect 636 -250 642 -246
rect 646 -247 650 -245
rect 694 -246 698 -235
rect 658 -247 698 -246
rect 658 -249 682 -247
rect 684 -249 698 -247
rect 658 -250 698 -249
rect 593 -257 594 -255
rect 596 -257 597 -255
rect 593 -259 597 -257
rect 602 -253 608 -252
rect 602 -255 604 -253
rect 606 -255 608 -253
rect 638 -254 662 -250
rect 681 -254 685 -250
rect 736 -215 746 -214
rect 736 -217 742 -215
rect 744 -217 746 -215
rect 736 -218 746 -217
rect 751 -215 772 -214
rect 751 -217 752 -215
rect 754 -216 772 -215
rect 774 -216 776 -214
rect 781 -215 785 -213
rect 754 -217 776 -216
rect 736 -222 740 -218
rect 720 -226 740 -222
rect 720 -229 724 -226
rect 718 -231 724 -229
rect 718 -233 719 -231
rect 721 -233 724 -231
rect 718 -235 724 -233
rect 720 -246 724 -235
rect 728 -231 732 -229
rect 751 -222 755 -217
rect 849 -215 869 -214
rect 849 -217 851 -215
rect 853 -217 869 -215
rect 849 -218 869 -217
rect 751 -224 752 -222
rect 754 -224 755 -222
rect 751 -226 755 -224
rect 760 -222 775 -221
rect 760 -224 762 -222
rect 764 -223 775 -222
rect 764 -224 789 -223
rect 760 -225 785 -224
rect 771 -226 785 -225
rect 787 -226 789 -224
rect 771 -227 789 -226
rect 728 -233 729 -231
rect 731 -233 732 -231
rect 728 -238 732 -233
rect 771 -238 775 -227
rect 768 -242 775 -238
rect 778 -234 782 -232
rect 778 -236 779 -234
rect 781 -236 782 -234
rect 768 -243 772 -242
rect 768 -245 769 -243
rect 771 -245 772 -243
rect 720 -247 760 -246
rect 768 -247 772 -245
rect 778 -246 782 -236
rect 811 -222 829 -221
rect 811 -224 813 -222
rect 815 -224 829 -222
rect 811 -225 829 -224
rect 825 -231 829 -225
rect 825 -233 826 -231
rect 828 -233 829 -231
rect 804 -238 810 -237
rect 720 -249 734 -247
rect 736 -249 760 -247
rect 720 -250 760 -249
rect 776 -250 782 -246
rect 733 -254 737 -250
rect 756 -254 780 -250
rect 825 -246 829 -233
rect 814 -250 829 -246
rect 814 -254 818 -250
rect 832 -254 833 -243
rect 865 -222 869 -218
rect 880 -221 881 -219
rect 865 -226 877 -222
rect 873 -231 877 -226
rect 873 -233 874 -231
rect 876 -233 877 -231
rect 873 -245 877 -233
rect 860 -248 877 -245
rect 860 -250 861 -248
rect 863 -249 877 -248
rect 863 -250 864 -249
rect 602 -264 608 -255
rect 668 -255 674 -254
rect 668 -257 670 -255
rect 672 -257 674 -255
rect 633 -262 639 -261
rect 633 -264 635 -262
rect 637 -264 639 -262
rect 668 -262 674 -257
rect 681 -256 682 -254
rect 684 -256 685 -254
rect 681 -258 685 -256
rect 690 -255 696 -254
rect 690 -257 692 -255
rect 694 -257 696 -255
rect 668 -264 670 -262
rect 672 -264 674 -262
rect 690 -262 696 -257
rect 690 -264 692 -262
rect 694 -264 696 -262
rect 722 -255 728 -254
rect 722 -257 724 -255
rect 726 -257 728 -255
rect 722 -262 728 -257
rect 733 -256 734 -254
rect 736 -256 737 -254
rect 733 -258 737 -256
rect 744 -255 750 -254
rect 744 -257 746 -255
rect 748 -257 750 -255
rect 722 -264 724 -262
rect 726 -264 728 -262
rect 744 -262 750 -257
rect 801 -255 818 -254
rect 801 -257 803 -255
rect 805 -257 818 -255
rect 801 -258 818 -257
rect 849 -255 855 -254
rect 849 -257 851 -255
rect 853 -257 855 -255
rect 744 -264 746 -262
rect 748 -264 750 -262
rect 779 -262 785 -261
rect 779 -264 781 -262
rect 783 -264 785 -262
rect 820 -262 826 -261
rect 820 -264 822 -262
rect 824 -264 826 -262
rect 849 -264 855 -257
rect 860 -255 864 -250
rect 900 -215 904 -213
rect 909 -214 934 -213
rect 1018 -214 1043 -213
rect 909 -216 911 -214
rect 913 -215 934 -214
rect 913 -216 931 -215
rect 909 -217 931 -216
rect 933 -217 934 -215
rect 910 -222 925 -221
rect 910 -223 921 -222
rect 896 -224 921 -223
rect 923 -224 925 -222
rect 896 -226 898 -224
rect 900 -225 925 -224
rect 930 -222 934 -217
rect 939 -215 949 -214
rect 939 -217 941 -215
rect 943 -217 949 -215
rect 939 -218 949 -217
rect 930 -224 931 -222
rect 933 -224 934 -222
rect 900 -226 914 -225
rect 930 -226 934 -224
rect 896 -227 914 -226
rect 903 -234 907 -232
rect 903 -236 904 -234
rect 906 -236 907 -234
rect 903 -246 907 -236
rect 910 -238 914 -227
rect 945 -222 949 -218
rect 945 -226 965 -222
rect 961 -229 965 -226
rect 953 -231 957 -229
rect 953 -233 954 -231
rect 956 -233 957 -231
rect 953 -238 957 -233
rect 961 -231 967 -229
rect 961 -233 964 -231
rect 966 -233 967 -231
rect 961 -235 967 -233
rect 910 -242 917 -238
rect 913 -243 917 -242
rect 913 -245 914 -243
rect 916 -245 917 -243
rect 903 -250 909 -246
rect 913 -247 917 -245
rect 961 -246 965 -235
rect 925 -247 965 -246
rect 925 -249 949 -247
rect 951 -249 965 -247
rect 925 -250 965 -249
rect 860 -257 861 -255
rect 863 -257 864 -255
rect 860 -259 864 -257
rect 869 -253 875 -252
rect 869 -255 871 -253
rect 873 -255 875 -253
rect 905 -254 929 -250
rect 948 -254 952 -250
rect 1003 -215 1013 -214
rect 1003 -217 1009 -215
rect 1011 -217 1013 -215
rect 1003 -218 1013 -217
rect 1018 -215 1039 -214
rect 1018 -217 1019 -215
rect 1021 -216 1039 -215
rect 1041 -216 1043 -214
rect 1048 -215 1052 -213
rect 1021 -217 1043 -216
rect 1003 -222 1007 -218
rect 987 -226 1007 -222
rect 987 -229 991 -226
rect 985 -231 991 -229
rect 985 -233 986 -231
rect 988 -233 991 -231
rect 985 -235 991 -233
rect 987 -246 991 -235
rect 995 -231 999 -229
rect 1018 -222 1022 -217
rect 1116 -215 1136 -214
rect 1116 -217 1118 -215
rect 1120 -217 1136 -215
rect 1116 -218 1136 -217
rect 1018 -224 1019 -222
rect 1021 -224 1022 -222
rect 1018 -226 1022 -224
rect 1027 -222 1042 -221
rect 1027 -224 1029 -222
rect 1031 -223 1042 -222
rect 1031 -224 1056 -223
rect 1027 -225 1052 -224
rect 1038 -226 1052 -225
rect 1054 -226 1056 -224
rect 1038 -227 1056 -226
rect 995 -233 996 -231
rect 998 -233 999 -231
rect 995 -238 999 -233
rect 1038 -238 1042 -227
rect 1035 -242 1042 -238
rect 1045 -234 1049 -232
rect 1045 -236 1046 -234
rect 1048 -236 1049 -234
rect 1035 -243 1039 -242
rect 1035 -245 1036 -243
rect 1038 -245 1039 -243
rect 987 -247 1027 -246
rect 1035 -247 1039 -245
rect 1045 -246 1049 -236
rect 1078 -222 1096 -221
rect 1078 -224 1080 -222
rect 1082 -224 1096 -222
rect 1078 -225 1096 -224
rect 1092 -231 1096 -225
rect 1092 -233 1093 -231
rect 1095 -233 1096 -231
rect 1071 -238 1077 -237
rect 987 -249 1001 -247
rect 1003 -249 1027 -247
rect 987 -250 1027 -249
rect 1043 -250 1049 -246
rect 1000 -254 1004 -250
rect 1023 -254 1047 -250
rect 1092 -246 1096 -233
rect 1081 -250 1096 -246
rect 1081 -254 1085 -250
rect 1099 -254 1100 -243
rect 1132 -222 1136 -218
rect 1147 -221 1148 -219
rect 1132 -226 1144 -222
rect 1140 -231 1144 -226
rect 1140 -233 1141 -231
rect 1143 -233 1144 -231
rect 1140 -245 1144 -233
rect 1127 -248 1144 -245
rect 1127 -250 1128 -248
rect 1130 -249 1144 -248
rect 1130 -250 1131 -249
rect 869 -264 875 -255
rect 935 -255 941 -254
rect 935 -257 937 -255
rect 939 -257 941 -255
rect 900 -262 906 -261
rect 900 -264 902 -262
rect 904 -264 906 -262
rect 935 -262 941 -257
rect 948 -256 949 -254
rect 951 -256 952 -254
rect 948 -258 952 -256
rect 957 -255 963 -254
rect 957 -257 959 -255
rect 961 -257 963 -255
rect 935 -264 937 -262
rect 939 -264 941 -262
rect 957 -262 963 -257
rect 957 -264 959 -262
rect 961 -264 963 -262
rect 989 -255 995 -254
rect 989 -257 991 -255
rect 993 -257 995 -255
rect 989 -262 995 -257
rect 1000 -256 1001 -254
rect 1003 -256 1004 -254
rect 1000 -258 1004 -256
rect 1011 -255 1017 -254
rect 1011 -257 1013 -255
rect 1015 -257 1017 -255
rect 989 -264 991 -262
rect 993 -264 995 -262
rect 1011 -262 1017 -257
rect 1068 -255 1085 -254
rect 1068 -257 1070 -255
rect 1072 -257 1085 -255
rect 1068 -258 1085 -257
rect 1116 -255 1122 -254
rect 1116 -257 1118 -255
rect 1120 -257 1122 -255
rect 1011 -264 1013 -262
rect 1015 -264 1017 -262
rect 1046 -262 1052 -261
rect 1046 -264 1048 -262
rect 1050 -264 1052 -262
rect 1087 -262 1093 -261
rect 1087 -264 1089 -262
rect 1091 -264 1093 -262
rect 1116 -264 1122 -257
rect 1127 -255 1131 -250
rect 1167 -215 1171 -213
rect 1176 -214 1201 -213
rect 1285 -214 1310 -213
rect 1176 -216 1178 -214
rect 1180 -215 1201 -214
rect 1180 -216 1198 -215
rect 1176 -217 1198 -216
rect 1200 -217 1201 -215
rect 1177 -222 1192 -221
rect 1177 -223 1188 -222
rect 1163 -224 1188 -223
rect 1190 -224 1192 -222
rect 1163 -226 1165 -224
rect 1167 -225 1192 -224
rect 1197 -222 1201 -217
rect 1206 -215 1216 -214
rect 1206 -217 1208 -215
rect 1210 -217 1216 -215
rect 1206 -218 1216 -217
rect 1197 -224 1198 -222
rect 1200 -224 1201 -222
rect 1167 -226 1181 -225
rect 1197 -226 1201 -224
rect 1163 -227 1181 -226
rect 1170 -234 1174 -232
rect 1170 -236 1171 -234
rect 1173 -236 1174 -234
rect 1170 -246 1174 -236
rect 1177 -238 1181 -227
rect 1212 -222 1216 -218
rect 1212 -226 1232 -222
rect 1228 -229 1232 -226
rect 1220 -231 1224 -229
rect 1220 -233 1221 -231
rect 1223 -233 1224 -231
rect 1220 -238 1224 -233
rect 1228 -231 1234 -229
rect 1228 -233 1231 -231
rect 1233 -233 1234 -231
rect 1228 -235 1234 -233
rect 1177 -242 1184 -238
rect 1180 -243 1184 -242
rect 1180 -245 1181 -243
rect 1183 -245 1184 -243
rect 1170 -250 1176 -246
rect 1180 -247 1184 -245
rect 1228 -246 1232 -235
rect 1192 -247 1232 -246
rect 1192 -249 1216 -247
rect 1218 -249 1232 -247
rect 1192 -250 1232 -249
rect 1127 -257 1128 -255
rect 1130 -257 1131 -255
rect 1127 -259 1131 -257
rect 1136 -253 1142 -252
rect 1136 -255 1138 -253
rect 1140 -255 1142 -253
rect 1172 -254 1196 -250
rect 1215 -254 1219 -250
rect 1270 -215 1280 -214
rect 1270 -217 1276 -215
rect 1278 -217 1280 -215
rect 1270 -218 1280 -217
rect 1285 -215 1306 -214
rect 1285 -217 1286 -215
rect 1288 -216 1306 -215
rect 1308 -216 1310 -214
rect 1315 -215 1319 -213
rect 1288 -217 1310 -216
rect 1270 -222 1274 -218
rect 1254 -226 1274 -222
rect 1254 -229 1258 -226
rect 1252 -231 1258 -229
rect 1252 -233 1253 -231
rect 1255 -233 1258 -231
rect 1252 -235 1258 -233
rect 1254 -246 1258 -235
rect 1262 -231 1266 -229
rect 1285 -222 1289 -217
rect 1383 -215 1403 -214
rect 1383 -217 1385 -215
rect 1387 -217 1403 -215
rect 1383 -218 1403 -217
rect 1285 -224 1286 -222
rect 1288 -224 1289 -222
rect 1285 -226 1289 -224
rect 1294 -222 1309 -221
rect 1294 -224 1296 -222
rect 1298 -223 1309 -222
rect 1298 -224 1323 -223
rect 1294 -225 1319 -224
rect 1305 -226 1319 -225
rect 1321 -226 1323 -224
rect 1305 -227 1323 -226
rect 1262 -233 1263 -231
rect 1265 -233 1266 -231
rect 1262 -238 1266 -233
rect 1305 -238 1309 -227
rect 1302 -242 1309 -238
rect 1312 -234 1316 -232
rect 1312 -236 1313 -234
rect 1315 -236 1316 -234
rect 1302 -243 1306 -242
rect 1302 -245 1303 -243
rect 1305 -245 1306 -243
rect 1254 -247 1294 -246
rect 1302 -247 1306 -245
rect 1312 -246 1316 -236
rect 1345 -222 1363 -221
rect 1345 -224 1347 -222
rect 1349 -224 1363 -222
rect 1345 -225 1363 -224
rect 1359 -231 1363 -225
rect 1359 -233 1360 -231
rect 1362 -233 1363 -231
rect 1338 -238 1344 -237
rect 1254 -249 1268 -247
rect 1270 -249 1294 -247
rect 1254 -250 1294 -249
rect 1310 -250 1316 -246
rect 1267 -254 1271 -250
rect 1290 -254 1314 -250
rect 1359 -246 1363 -233
rect 1348 -250 1363 -246
rect 1348 -254 1352 -250
rect 1366 -254 1367 -243
rect 1399 -222 1403 -218
rect 1414 -221 1415 -219
rect 1399 -226 1411 -222
rect 1407 -231 1411 -226
rect 1407 -233 1408 -231
rect 1410 -233 1411 -231
rect 1407 -245 1411 -233
rect 1394 -248 1411 -245
rect 1394 -250 1395 -248
rect 1397 -249 1411 -248
rect 1397 -250 1398 -249
rect 1136 -264 1142 -255
rect 1202 -255 1208 -254
rect 1202 -257 1204 -255
rect 1206 -257 1208 -255
rect 1167 -262 1173 -261
rect 1167 -264 1169 -262
rect 1171 -264 1173 -262
rect 1202 -262 1208 -257
rect 1215 -256 1216 -254
rect 1218 -256 1219 -254
rect 1215 -258 1219 -256
rect 1224 -255 1230 -254
rect 1224 -257 1226 -255
rect 1228 -257 1230 -255
rect 1202 -264 1204 -262
rect 1206 -264 1208 -262
rect 1224 -262 1230 -257
rect 1224 -264 1226 -262
rect 1228 -264 1230 -262
rect 1256 -255 1262 -254
rect 1256 -257 1258 -255
rect 1260 -257 1262 -255
rect 1256 -262 1262 -257
rect 1267 -256 1268 -254
rect 1270 -256 1271 -254
rect 1267 -258 1271 -256
rect 1278 -255 1284 -254
rect 1278 -257 1280 -255
rect 1282 -257 1284 -255
rect 1256 -264 1258 -262
rect 1260 -264 1262 -262
rect 1278 -262 1284 -257
rect 1335 -255 1352 -254
rect 1335 -257 1337 -255
rect 1339 -257 1352 -255
rect 1335 -258 1352 -257
rect 1383 -255 1389 -254
rect 1383 -257 1385 -255
rect 1387 -257 1389 -255
rect 1278 -264 1280 -262
rect 1282 -264 1284 -262
rect 1313 -262 1319 -261
rect 1313 -264 1315 -262
rect 1317 -264 1319 -262
rect 1354 -262 1360 -261
rect 1354 -264 1356 -262
rect 1358 -264 1360 -262
rect 1383 -264 1389 -257
rect 1394 -255 1398 -250
rect 1434 -215 1438 -213
rect 1443 -214 1468 -213
rect 1552 -214 1577 -213
rect 1443 -216 1445 -214
rect 1447 -215 1468 -214
rect 1447 -216 1465 -215
rect 1443 -217 1465 -216
rect 1467 -217 1468 -215
rect 1444 -222 1459 -221
rect 1444 -223 1455 -222
rect 1430 -224 1455 -223
rect 1457 -224 1459 -222
rect 1430 -226 1432 -224
rect 1434 -225 1459 -224
rect 1464 -222 1468 -217
rect 1473 -215 1483 -214
rect 1473 -217 1475 -215
rect 1477 -217 1483 -215
rect 1473 -218 1483 -217
rect 1464 -224 1465 -222
rect 1467 -224 1468 -222
rect 1434 -226 1448 -225
rect 1464 -226 1468 -224
rect 1430 -227 1448 -226
rect 1437 -234 1441 -232
rect 1437 -236 1438 -234
rect 1440 -236 1441 -234
rect 1437 -246 1441 -236
rect 1444 -238 1448 -227
rect 1479 -222 1483 -218
rect 1479 -226 1499 -222
rect 1495 -229 1499 -226
rect 1487 -231 1491 -229
rect 1487 -233 1488 -231
rect 1490 -233 1491 -231
rect 1487 -238 1491 -233
rect 1495 -231 1501 -229
rect 1495 -233 1498 -231
rect 1500 -233 1501 -231
rect 1495 -235 1501 -233
rect 1444 -242 1451 -238
rect 1447 -243 1451 -242
rect 1447 -245 1448 -243
rect 1450 -245 1451 -243
rect 1437 -250 1443 -246
rect 1447 -247 1451 -245
rect 1495 -246 1499 -235
rect 1459 -247 1499 -246
rect 1459 -249 1483 -247
rect 1485 -249 1499 -247
rect 1459 -250 1499 -249
rect 1394 -257 1395 -255
rect 1397 -257 1398 -255
rect 1394 -259 1398 -257
rect 1403 -253 1409 -252
rect 1403 -255 1405 -253
rect 1407 -255 1409 -253
rect 1439 -254 1463 -250
rect 1482 -254 1486 -250
rect 1537 -215 1547 -214
rect 1537 -217 1543 -215
rect 1545 -217 1547 -215
rect 1537 -218 1547 -217
rect 1552 -215 1573 -214
rect 1552 -217 1553 -215
rect 1555 -216 1573 -215
rect 1575 -216 1577 -214
rect 1582 -215 1586 -213
rect 1555 -217 1577 -216
rect 1537 -222 1541 -218
rect 1521 -226 1541 -222
rect 1521 -229 1525 -226
rect 1519 -231 1525 -229
rect 1519 -233 1520 -231
rect 1522 -233 1525 -231
rect 1519 -235 1525 -233
rect 1521 -246 1525 -235
rect 1529 -231 1533 -229
rect 1552 -222 1556 -217
rect 1650 -215 1670 -214
rect 1650 -217 1652 -215
rect 1654 -217 1670 -215
rect 1650 -218 1670 -217
rect 1552 -224 1553 -222
rect 1555 -224 1556 -222
rect 1552 -226 1556 -224
rect 1561 -222 1576 -221
rect 1561 -224 1563 -222
rect 1565 -223 1576 -222
rect 1565 -224 1590 -223
rect 1561 -225 1586 -224
rect 1572 -226 1586 -225
rect 1588 -226 1590 -224
rect 1572 -227 1590 -226
rect 1529 -233 1530 -231
rect 1532 -233 1533 -231
rect 1529 -238 1533 -233
rect 1572 -238 1576 -227
rect 1569 -242 1576 -238
rect 1579 -234 1583 -232
rect 1579 -236 1580 -234
rect 1582 -236 1583 -234
rect 1569 -243 1573 -242
rect 1569 -245 1570 -243
rect 1572 -245 1573 -243
rect 1521 -247 1561 -246
rect 1569 -247 1573 -245
rect 1579 -246 1583 -236
rect 1612 -222 1630 -221
rect 1612 -224 1614 -222
rect 1616 -224 1630 -222
rect 1612 -225 1630 -224
rect 1626 -231 1630 -225
rect 1626 -233 1627 -231
rect 1629 -233 1630 -231
rect 1605 -238 1611 -237
rect 1521 -249 1535 -247
rect 1537 -249 1561 -247
rect 1521 -250 1561 -249
rect 1577 -250 1583 -246
rect 1534 -254 1538 -250
rect 1557 -254 1581 -250
rect 1626 -246 1630 -233
rect 1615 -250 1630 -246
rect 1615 -254 1619 -250
rect 1633 -254 1634 -243
rect 1666 -222 1670 -218
rect 1681 -221 1682 -219
rect 1666 -226 1678 -222
rect 1674 -231 1678 -226
rect 1674 -233 1675 -231
rect 1677 -233 1678 -231
rect 1674 -245 1678 -233
rect 1661 -248 1678 -245
rect 1661 -250 1662 -248
rect 1664 -249 1678 -248
rect 1664 -250 1665 -249
rect 1403 -264 1409 -255
rect 1469 -255 1475 -254
rect 1469 -257 1471 -255
rect 1473 -257 1475 -255
rect 1434 -262 1440 -261
rect 1434 -264 1436 -262
rect 1438 -264 1440 -262
rect 1469 -262 1475 -257
rect 1482 -256 1483 -254
rect 1485 -256 1486 -254
rect 1482 -258 1486 -256
rect 1491 -255 1497 -254
rect 1491 -257 1493 -255
rect 1495 -257 1497 -255
rect 1469 -264 1471 -262
rect 1473 -264 1475 -262
rect 1491 -262 1497 -257
rect 1491 -264 1493 -262
rect 1495 -264 1497 -262
rect 1523 -255 1529 -254
rect 1523 -257 1525 -255
rect 1527 -257 1529 -255
rect 1523 -262 1529 -257
rect 1534 -256 1535 -254
rect 1537 -256 1538 -254
rect 1534 -258 1538 -256
rect 1545 -255 1551 -254
rect 1545 -257 1547 -255
rect 1549 -257 1551 -255
rect 1523 -264 1525 -262
rect 1527 -264 1529 -262
rect 1545 -262 1551 -257
rect 1602 -255 1619 -254
rect 1602 -257 1604 -255
rect 1606 -257 1619 -255
rect 1602 -258 1619 -257
rect 1650 -255 1656 -254
rect 1650 -257 1652 -255
rect 1654 -257 1656 -255
rect 1545 -264 1547 -262
rect 1549 -264 1551 -262
rect 1580 -262 1586 -261
rect 1580 -264 1582 -262
rect 1584 -264 1586 -262
rect 1621 -262 1627 -261
rect 1621 -264 1623 -262
rect 1625 -264 1627 -262
rect 1650 -264 1656 -257
rect 1661 -255 1665 -250
rect 1701 -215 1705 -213
rect 1710 -214 1735 -213
rect 1819 -214 1844 -213
rect 1710 -216 1712 -214
rect 1714 -215 1735 -214
rect 1714 -216 1732 -215
rect 1710 -217 1732 -216
rect 1734 -217 1735 -215
rect 1711 -222 1726 -221
rect 1711 -223 1722 -222
rect 1697 -224 1722 -223
rect 1724 -224 1726 -222
rect 1697 -226 1699 -224
rect 1701 -225 1726 -224
rect 1731 -222 1735 -217
rect 1740 -215 1750 -214
rect 1740 -217 1742 -215
rect 1744 -217 1750 -215
rect 1740 -218 1750 -217
rect 1731 -224 1732 -222
rect 1734 -224 1735 -222
rect 1701 -226 1715 -225
rect 1731 -226 1735 -224
rect 1697 -227 1715 -226
rect 1704 -234 1708 -232
rect 1704 -236 1705 -234
rect 1707 -236 1708 -234
rect 1704 -246 1708 -236
rect 1711 -238 1715 -227
rect 1746 -222 1750 -218
rect 1746 -226 1766 -222
rect 1762 -229 1766 -226
rect 1754 -231 1758 -229
rect 1754 -233 1755 -231
rect 1757 -233 1758 -231
rect 1754 -238 1758 -233
rect 1762 -231 1768 -229
rect 1762 -233 1765 -231
rect 1767 -233 1768 -231
rect 1762 -235 1768 -233
rect 1711 -242 1718 -238
rect 1714 -243 1718 -242
rect 1714 -245 1715 -243
rect 1717 -245 1718 -243
rect 1704 -250 1710 -246
rect 1714 -247 1718 -245
rect 1762 -246 1766 -235
rect 1726 -247 1766 -246
rect 1726 -249 1750 -247
rect 1752 -249 1766 -247
rect 1726 -250 1766 -249
rect 1661 -257 1662 -255
rect 1664 -257 1665 -255
rect 1661 -259 1665 -257
rect 1670 -253 1676 -252
rect 1670 -255 1672 -253
rect 1674 -255 1676 -253
rect 1706 -254 1730 -250
rect 1749 -254 1753 -250
rect 1804 -215 1814 -214
rect 1804 -217 1810 -215
rect 1812 -217 1814 -215
rect 1804 -218 1814 -217
rect 1819 -215 1840 -214
rect 1819 -217 1820 -215
rect 1822 -216 1840 -215
rect 1842 -216 1844 -214
rect 1849 -215 1853 -213
rect 1822 -217 1844 -216
rect 1926 -214 1932 -208
rect 1987 -211 1991 -208
rect 2043 -210 2045 -208
rect 2047 -210 2049 -208
rect 2043 -211 2049 -210
rect 2077 -210 2079 -208
rect 2081 -210 2083 -208
rect 2077 -211 2083 -210
rect 2135 -211 2139 -208
rect 1987 -213 1988 -211
rect 1990 -213 1991 -211
rect 2135 -213 2136 -211
rect 2138 -213 2139 -211
rect 2155 -209 2161 -208
rect 2155 -211 2157 -209
rect 2159 -211 2161 -209
rect 2155 -212 2161 -211
rect 2174 -209 2180 -208
rect 2174 -211 2176 -209
rect 2178 -211 2180 -209
rect 2174 -212 2180 -211
rect 1926 -216 1928 -214
rect 1930 -216 1932 -214
rect 1926 -217 1932 -216
rect 1939 -217 1943 -215
rect 1804 -222 1808 -218
rect 1788 -226 1808 -222
rect 1788 -229 1792 -226
rect 1786 -231 1792 -229
rect 1786 -233 1787 -231
rect 1789 -233 1792 -231
rect 1786 -235 1792 -233
rect 1788 -246 1792 -235
rect 1796 -231 1800 -229
rect 1819 -222 1823 -217
rect 1939 -219 1940 -217
rect 1942 -219 1943 -217
rect 1819 -224 1820 -222
rect 1822 -224 1823 -222
rect 1819 -226 1823 -224
rect 1828 -222 1843 -221
rect 1828 -224 1830 -222
rect 1832 -223 1843 -222
rect 1832 -224 1857 -223
rect 1828 -225 1853 -224
rect 1839 -226 1853 -225
rect 1855 -226 1857 -224
rect 1839 -227 1857 -226
rect 1796 -233 1797 -231
rect 1799 -233 1800 -231
rect 1796 -238 1800 -233
rect 1839 -238 1843 -227
rect 1836 -242 1843 -238
rect 1846 -234 1850 -232
rect 1846 -236 1847 -234
rect 1849 -236 1850 -234
rect 1836 -243 1840 -242
rect 1836 -245 1837 -243
rect 1839 -245 1840 -243
rect 1788 -247 1828 -246
rect 1836 -247 1840 -245
rect 1846 -246 1850 -236
rect 1879 -222 1897 -221
rect 1879 -224 1881 -222
rect 1883 -224 1897 -222
rect 1879 -225 1897 -224
rect 1893 -231 1897 -225
rect 1893 -233 1894 -231
rect 1896 -233 1897 -231
rect 1872 -238 1878 -237
rect 1788 -249 1802 -247
rect 1804 -249 1828 -247
rect 1788 -250 1828 -249
rect 1844 -250 1850 -246
rect 1801 -254 1805 -250
rect 1824 -254 1848 -250
rect 1893 -246 1897 -233
rect 1882 -250 1897 -246
rect 1882 -254 1886 -250
rect 1900 -254 1901 -243
rect 1913 -222 1917 -220
rect 1913 -224 1914 -222
rect 1916 -224 1917 -222
rect 1913 -230 1917 -224
rect 1939 -222 1943 -219
rect 1939 -226 1963 -222
rect 1913 -234 1924 -230
rect 1670 -264 1676 -255
rect 1736 -255 1742 -254
rect 1736 -257 1738 -255
rect 1740 -257 1742 -255
rect 1701 -262 1707 -261
rect 1701 -264 1703 -262
rect 1705 -264 1707 -262
rect 1736 -262 1742 -257
rect 1749 -256 1750 -254
rect 1752 -256 1753 -254
rect 1749 -258 1753 -256
rect 1758 -255 1764 -254
rect 1758 -257 1760 -255
rect 1762 -257 1764 -255
rect 1736 -264 1738 -262
rect 1740 -264 1742 -262
rect 1758 -262 1764 -257
rect 1758 -264 1760 -262
rect 1762 -264 1764 -262
rect 1790 -255 1796 -254
rect 1790 -257 1792 -255
rect 1794 -257 1796 -255
rect 1790 -262 1796 -257
rect 1801 -256 1802 -254
rect 1804 -256 1805 -254
rect 1801 -258 1805 -256
rect 1812 -255 1818 -254
rect 1812 -257 1814 -255
rect 1816 -257 1818 -255
rect 1790 -264 1792 -262
rect 1794 -264 1796 -262
rect 1812 -262 1818 -257
rect 1869 -255 1886 -254
rect 1869 -257 1871 -255
rect 1873 -257 1886 -255
rect 1869 -258 1886 -257
rect 1920 -240 1924 -234
rect 1959 -230 1963 -226
rect 1939 -231 1955 -230
rect 1939 -233 1951 -231
rect 1953 -233 1955 -231
rect 1939 -234 1955 -233
rect 1959 -232 1964 -230
rect 1959 -234 1961 -232
rect 1963 -234 1964 -232
rect 1939 -240 1943 -234
rect 1959 -236 1964 -234
rect 1959 -238 1963 -236
rect 1920 -241 1943 -240
rect 1920 -243 1922 -241
rect 1924 -243 1943 -241
rect 1920 -244 1943 -243
rect 1931 -255 1935 -253
rect 1931 -257 1932 -255
rect 1934 -257 1935 -255
rect 1812 -264 1814 -262
rect 1816 -264 1818 -262
rect 1847 -262 1853 -261
rect 1847 -264 1849 -262
rect 1851 -264 1853 -262
rect 1888 -262 1894 -261
rect 1888 -264 1890 -262
rect 1892 -264 1894 -262
rect 1931 -262 1935 -257
rect 1939 -255 1943 -244
rect 1947 -241 1963 -238
rect 1947 -243 1948 -241
rect 1950 -242 1963 -241
rect 1950 -243 1951 -242
rect 1947 -248 1951 -243
rect 1947 -250 1948 -248
rect 1950 -250 1951 -248
rect 1947 -252 1951 -250
rect 1987 -215 1991 -213
rect 1996 -214 2021 -213
rect 2105 -214 2130 -213
rect 1996 -216 1998 -214
rect 2000 -215 2021 -214
rect 2000 -216 2018 -215
rect 1996 -217 2018 -216
rect 2020 -217 2021 -215
rect 1997 -222 2012 -221
rect 1997 -223 2008 -222
rect 1983 -224 2008 -223
rect 2010 -224 2012 -222
rect 1983 -226 1985 -224
rect 1987 -225 2012 -224
rect 2017 -222 2021 -217
rect 2026 -215 2036 -214
rect 2026 -217 2028 -215
rect 2030 -217 2036 -215
rect 2026 -218 2036 -217
rect 2017 -224 2018 -222
rect 2020 -224 2021 -222
rect 1987 -226 2001 -225
rect 2017 -226 2021 -224
rect 1983 -227 2001 -226
rect 1990 -234 1994 -232
rect 1990 -236 1991 -234
rect 1993 -236 1994 -234
rect 1990 -246 1994 -236
rect 1997 -238 2001 -227
rect 2032 -222 2036 -218
rect 2032 -226 2052 -222
rect 2048 -229 2052 -226
rect 2040 -231 2044 -229
rect 2040 -233 2041 -231
rect 2043 -233 2044 -231
rect 2040 -238 2044 -233
rect 2048 -231 2054 -229
rect 2048 -233 2051 -231
rect 2053 -233 2054 -231
rect 2048 -235 2054 -233
rect 1997 -242 2004 -238
rect 2000 -243 2004 -242
rect 2000 -245 2001 -243
rect 2003 -245 2004 -243
rect 1990 -250 1996 -246
rect 2000 -247 2004 -245
rect 2048 -246 2052 -235
rect 2012 -247 2052 -246
rect 2012 -249 2036 -247
rect 2038 -249 2052 -247
rect 2012 -250 2052 -249
rect 1992 -254 2016 -250
rect 2035 -254 2039 -250
rect 2090 -215 2100 -214
rect 2090 -217 2096 -215
rect 2098 -217 2100 -215
rect 2090 -218 2100 -217
rect 2105 -215 2126 -214
rect 2105 -217 2106 -215
rect 2108 -216 2126 -215
rect 2128 -216 2130 -214
rect 2135 -215 2139 -213
rect 2108 -217 2130 -216
rect 2199 -216 2205 -215
rect 2090 -222 2094 -218
rect 2074 -226 2094 -222
rect 2074 -229 2078 -226
rect 2072 -231 2078 -229
rect 2072 -233 2073 -231
rect 2075 -233 2078 -231
rect 2072 -235 2078 -233
rect 2074 -246 2078 -235
rect 2082 -231 2086 -229
rect 2105 -222 2109 -217
rect 2105 -224 2106 -222
rect 2108 -224 2109 -222
rect 2105 -226 2109 -224
rect 2114 -222 2129 -221
rect 2114 -224 2116 -222
rect 2118 -223 2129 -222
rect 2118 -224 2143 -223
rect 2114 -225 2139 -224
rect 2125 -226 2139 -225
rect 2141 -226 2143 -224
rect 2125 -227 2143 -226
rect 2082 -233 2083 -231
rect 2085 -233 2086 -231
rect 2082 -238 2086 -233
rect 2125 -238 2129 -227
rect 2122 -242 2129 -238
rect 2132 -234 2136 -232
rect 2132 -236 2133 -234
rect 2135 -236 2136 -234
rect 2122 -243 2126 -242
rect 2122 -245 2123 -243
rect 2125 -245 2126 -243
rect 2074 -247 2114 -246
rect 2122 -247 2126 -245
rect 2132 -246 2136 -236
rect 2199 -218 2201 -216
rect 2203 -218 2205 -216
rect 2199 -219 2205 -218
rect 2209 -216 2215 -208
rect 2209 -218 2211 -216
rect 2213 -218 2215 -216
rect 2226 -214 2241 -213
rect 2226 -216 2228 -214
rect 2230 -216 2241 -214
rect 2226 -217 2241 -216
rect 2209 -219 2215 -218
rect 2165 -222 2183 -221
rect 2165 -224 2167 -222
rect 2169 -224 2183 -222
rect 2165 -225 2183 -224
rect 2179 -231 2183 -225
rect 2179 -233 2180 -231
rect 2182 -233 2183 -231
rect 2158 -238 2164 -237
rect 2074 -249 2088 -247
rect 2090 -249 2114 -247
rect 2074 -250 2114 -249
rect 2130 -250 2136 -246
rect 2087 -254 2091 -250
rect 2110 -254 2134 -250
rect 2179 -246 2183 -233
rect 2168 -250 2183 -246
rect 2168 -254 2172 -250
rect 2186 -254 2187 -243
rect 2199 -239 2203 -219
rect 2237 -222 2241 -217
rect 2244 -214 2248 -208
rect 2244 -216 2245 -214
rect 2247 -216 2248 -214
rect 2244 -218 2248 -216
rect 2223 -225 2234 -223
rect 2223 -227 2231 -225
rect 2233 -227 2234 -225
rect 2237 -224 2251 -222
rect 2237 -226 2252 -224
rect 2223 -229 2234 -227
rect 2247 -228 2249 -226
rect 2251 -228 2252 -226
rect 2223 -239 2227 -229
rect 2247 -230 2252 -228
rect 2199 -240 2227 -239
rect 2199 -242 2201 -240
rect 2203 -241 2227 -240
rect 2203 -242 2224 -241
rect 2199 -243 2224 -242
rect 2226 -243 2227 -241
rect 2243 -240 2244 -234
rect 2223 -245 2227 -243
rect 2022 -255 2028 -254
rect 1939 -256 1972 -255
rect 1939 -258 1968 -256
rect 1970 -258 1972 -256
rect 1939 -259 1972 -258
rect 2022 -257 2024 -255
rect 2026 -257 2028 -255
rect 1931 -264 1932 -262
rect 1934 -264 1935 -262
rect 1987 -262 1993 -261
rect 1987 -264 1989 -262
rect 1991 -264 1993 -262
rect 2022 -262 2028 -257
rect 2035 -256 2036 -254
rect 2038 -256 2039 -254
rect 2035 -258 2039 -256
rect 2044 -255 2050 -254
rect 2044 -257 2046 -255
rect 2048 -257 2050 -255
rect 2022 -264 2024 -262
rect 2026 -264 2028 -262
rect 2044 -262 2050 -257
rect 2044 -264 2046 -262
rect 2048 -264 2050 -262
rect 2076 -255 2082 -254
rect 2076 -257 2078 -255
rect 2080 -257 2082 -255
rect 2076 -262 2082 -257
rect 2087 -256 2088 -254
rect 2090 -256 2091 -254
rect 2087 -258 2091 -256
rect 2098 -255 2104 -254
rect 2098 -257 2100 -255
rect 2102 -257 2104 -255
rect 2076 -264 2078 -262
rect 2080 -264 2082 -262
rect 2098 -262 2104 -257
rect 2155 -255 2172 -254
rect 2155 -257 2157 -255
rect 2159 -257 2172 -255
rect 2155 -258 2172 -257
rect 2247 -247 2251 -230
rect 2235 -251 2251 -247
rect 2226 -252 2239 -251
rect 2226 -254 2228 -252
rect 2230 -254 2239 -252
rect 2267 -216 2273 -215
rect 2267 -218 2269 -216
rect 2271 -218 2273 -216
rect 2267 -219 2273 -218
rect 2277 -216 2283 -208
rect 2277 -218 2279 -216
rect 2281 -218 2283 -216
rect 2294 -214 2309 -213
rect 2294 -216 2296 -214
rect 2298 -216 2309 -214
rect 2294 -217 2309 -216
rect 2277 -219 2283 -218
rect 2267 -239 2271 -219
rect 2305 -222 2309 -217
rect 2312 -214 2316 -208
rect 2312 -216 2313 -214
rect 2315 -216 2316 -214
rect 2312 -218 2316 -216
rect 2291 -225 2302 -223
rect 2291 -227 2299 -225
rect 2301 -227 2302 -225
rect 2305 -224 2319 -222
rect 2305 -226 2320 -224
rect 2291 -229 2302 -227
rect 2315 -228 2317 -226
rect 2319 -228 2320 -226
rect 2291 -239 2295 -229
rect 2315 -230 2320 -228
rect 2267 -240 2295 -239
rect 2267 -242 2269 -240
rect 2271 -241 2295 -240
rect 2271 -242 2292 -241
rect 2267 -243 2292 -242
rect 2294 -243 2295 -241
rect 2311 -240 2312 -234
rect 2291 -245 2295 -243
rect 2226 -255 2239 -254
rect 2315 -247 2319 -230
rect 2303 -251 2319 -247
rect 2294 -252 2307 -251
rect 2294 -254 2296 -252
rect 2298 -254 2307 -252
rect 2294 -255 2307 -254
rect 2098 -264 2100 -262
rect 2102 -264 2104 -262
rect 2133 -262 2139 -261
rect 2133 -264 2135 -262
rect 2137 -264 2139 -262
rect 2174 -262 2180 -261
rect 2174 -264 2176 -262
rect 2178 -264 2180 -262
rect 2210 -262 2214 -260
rect 2210 -264 2211 -262
rect 2213 -264 2214 -262
rect 2243 -262 2249 -261
rect 2243 -264 2245 -262
rect 2247 -264 2249 -262
rect 2278 -262 2282 -260
rect 2278 -264 2279 -262
rect 2281 -264 2282 -262
rect 2311 -262 2317 -261
rect 2311 -264 2313 -262
rect 2315 -264 2317 -262
<< via1 >>
rect 2320 301 2322 303
rect 9 274 11 276
rect 41 268 43 270
rect 57 257 59 259
rect 81 263 83 265
rect 121 271 123 273
rect 139 263 141 265
rect 89 255 91 257
rect 170 263 172 265
rect 180 276 182 278
rect 210 271 212 273
rect 259 271 261 273
rect 211 255 213 257
rect 268 280 270 282
rect 268 263 270 265
rect 300 259 302 261
rect 324 257 326 259
rect 348 263 350 265
rect 388 271 390 273
rect 406 263 408 265
rect 356 255 358 257
rect 437 263 439 265
rect 447 276 449 278
rect 477 271 479 273
rect 526 271 528 273
rect 478 255 480 257
rect 535 280 537 282
rect 535 263 537 265
rect 567 259 569 261
rect 591 257 593 259
rect 615 263 617 265
rect 655 271 657 273
rect 673 263 675 265
rect 623 255 625 257
rect 704 263 706 265
rect 714 276 716 278
rect 744 271 746 273
rect 745 255 747 257
rect 802 280 804 282
rect 793 255 795 257
rect 802 263 804 265
rect 834 259 836 261
rect 858 257 860 259
rect 882 263 884 265
rect 922 271 924 273
rect 940 263 942 265
rect 890 255 892 257
rect 971 263 973 265
rect 981 276 983 278
rect 1011 271 1013 273
rect 1012 255 1014 257
rect 1069 280 1071 282
rect 1060 255 1062 257
rect 1069 263 1071 265
rect 1101 259 1103 261
rect 1125 257 1127 259
rect 1149 263 1151 265
rect 1189 271 1191 273
rect 1207 263 1209 265
rect 1157 255 1159 257
rect 1238 263 1240 265
rect 1248 276 1250 278
rect 1278 271 1280 273
rect 1279 255 1281 257
rect 1336 280 1338 282
rect 1327 252 1329 254
rect 1336 263 1338 265
rect 1368 259 1370 261
rect 1392 257 1394 259
rect 1416 263 1418 265
rect 1456 271 1458 273
rect 1474 263 1476 265
rect 1424 255 1426 257
rect 1505 263 1507 265
rect 1515 276 1517 278
rect 1545 271 1547 273
rect 1546 255 1548 257
rect 1603 280 1605 282
rect 1594 252 1596 254
rect 1603 263 1605 265
rect 1635 259 1637 261
rect 1659 257 1661 259
rect 1683 263 1685 265
rect 1723 271 1725 273
rect 1741 263 1743 265
rect 1691 255 1693 257
rect 1772 263 1774 265
rect 1782 276 1784 278
rect 1812 271 1814 273
rect 1861 271 1863 273
rect 1813 255 1815 257
rect 1870 280 1872 282
rect 1870 263 1872 265
rect 1902 259 1904 261
rect 1969 271 1971 273
rect 1925 254 1927 256
rect 2018 271 2020 273
rect 1977 255 1979 257
rect 2058 263 2060 265
rect 2068 276 2070 278
rect 2100 271 2102 273
rect 2099 255 2101 257
rect 2156 276 2158 278
rect 2147 255 2149 257
rect 2156 263 2158 265
rect 2188 259 2190 261
rect 2208 255 2210 257
rect 2236 271 2238 273
rect 2276 255 2278 257
rect 2300 272 2302 274
rect 216 234 218 236
rect 483 234 485 236
rect 750 234 752 236
rect 1017 234 1019 236
rect 1284 234 1286 236
rect 1551 234 1553 236
rect 1818 234 1820 236
rect 2276 231 2278 233
rect 2311 227 2313 229
rect 17 203 19 205
rect 41 191 43 193
rect 81 199 83 201
rect 49 183 51 185
rect 89 207 91 209
rect 139 199 141 201
rect 170 199 172 201
rect 134 191 136 193
rect 261 216 263 218
rect 211 207 213 209
rect 180 186 182 188
rect 228 194 230 196
rect 268 205 270 207
rect 268 186 270 188
rect 348 199 350 201
rect 316 183 318 185
rect 292 175 294 177
rect 356 207 358 209
rect 406 199 408 201
rect 437 199 439 201
rect 401 191 403 193
rect 528 216 530 218
rect 478 207 480 209
rect 447 186 449 188
rect 495 194 497 196
rect 535 205 537 207
rect 535 186 537 188
rect 615 199 617 201
rect 583 183 585 185
rect 559 175 561 177
rect 623 207 625 209
rect 673 199 675 201
rect 704 199 706 201
rect 668 191 670 193
rect 795 216 797 218
rect 745 207 747 209
rect 714 186 716 188
rect 762 194 764 196
rect 802 205 804 207
rect 802 186 804 188
rect 882 199 884 201
rect 850 183 852 185
rect 826 175 828 177
rect 890 207 892 209
rect 940 199 942 201
rect 971 199 973 201
rect 935 191 937 193
rect 1062 216 1064 218
rect 1012 207 1014 209
rect 981 186 983 188
rect 1029 194 1031 196
rect 1069 205 1071 207
rect 1069 186 1071 188
rect 1149 199 1151 201
rect 1117 183 1119 185
rect 1093 175 1095 177
rect 1157 207 1159 209
rect 1207 199 1209 201
rect 1238 199 1240 201
rect 1202 191 1204 193
rect 1329 216 1331 218
rect 1279 207 1281 209
rect 1248 186 1250 188
rect 1296 194 1298 196
rect 1336 205 1338 207
rect 1336 186 1338 188
rect 1416 199 1418 201
rect 1384 183 1386 185
rect 1360 175 1362 177
rect 1424 207 1426 209
rect 1474 199 1476 201
rect 1505 199 1507 201
rect 1469 191 1471 193
rect 1596 216 1598 218
rect 1546 207 1548 209
rect 1515 186 1517 188
rect 1563 194 1565 196
rect 1603 205 1605 207
rect 1603 186 1605 188
rect 1683 199 1685 201
rect 1651 183 1653 185
rect 1627 175 1629 177
rect 1691 207 1693 209
rect 1741 199 1743 201
rect 1772 199 1774 201
rect 1736 191 1738 193
rect 1863 216 1865 218
rect 1813 207 1815 209
rect 1782 186 1784 188
rect 1830 194 1832 196
rect 1870 205 1872 207
rect 1870 186 1872 188
rect 1925 208 1927 210
rect 1894 175 1896 177
rect 1969 191 1971 193
rect 1977 207 1979 209
rect 2058 199 2060 201
rect 2018 191 2020 193
rect 2149 216 2151 218
rect 2099 207 2101 209
rect 2068 186 2070 188
rect 2116 194 2118 196
rect 2156 205 2158 207
rect 2156 186 2158 188
rect 2210 207 2212 209
rect 2236 191 2238 193
rect 2180 175 2182 177
rect 2276 207 2278 209
rect 2300 192 2302 194
rect 2320 165 2322 167
rect 9 130 11 132
rect 41 127 43 129
rect 57 114 59 116
rect 81 119 83 121
rect 138 127 140 129
rect 140 119 142 121
rect 89 111 91 113
rect 170 119 172 121
rect 180 132 182 134
rect 228 127 230 129
rect 211 111 213 113
rect 268 136 270 138
rect 268 119 270 121
rect 300 115 302 117
rect 324 114 326 116
rect 348 119 350 121
rect 261 102 263 104
rect 405 127 407 129
rect 407 119 409 121
rect 356 111 358 113
rect 437 119 439 121
rect 447 132 449 134
rect 495 127 497 129
rect 478 111 480 113
rect 535 136 537 138
rect 535 119 537 121
rect 567 115 569 117
rect 591 114 593 116
rect 615 119 617 121
rect 528 102 530 104
rect 672 127 674 129
rect 674 119 676 121
rect 623 111 625 113
rect 704 119 706 121
rect 714 132 716 134
rect 762 127 764 129
rect 745 111 747 113
rect 802 136 804 138
rect 802 119 804 121
rect 834 115 836 117
rect 858 114 860 116
rect 882 119 884 121
rect 795 102 797 104
rect 939 127 941 129
rect 941 119 943 121
rect 890 111 892 113
rect 971 119 973 121
rect 981 132 983 134
rect 1029 127 1031 129
rect 1012 111 1014 113
rect 1069 136 1071 138
rect 1069 119 1071 121
rect 1101 115 1103 117
rect 1125 114 1127 116
rect 1149 119 1151 121
rect 1062 102 1064 104
rect 1206 127 1208 129
rect 1208 119 1210 121
rect 1157 111 1159 113
rect 1238 119 1240 121
rect 1248 132 1250 134
rect 1296 127 1298 129
rect 1279 111 1281 113
rect 1336 136 1338 138
rect 1336 119 1338 121
rect 1368 115 1370 117
rect 1392 114 1394 116
rect 1416 119 1418 121
rect 1329 102 1331 104
rect 1473 127 1475 129
rect 1475 119 1477 121
rect 1424 111 1426 113
rect 1505 119 1507 121
rect 1515 132 1517 134
rect 1563 127 1565 129
rect 1546 111 1548 113
rect 1603 136 1605 138
rect 1603 119 1605 121
rect 1635 115 1637 117
rect 1659 114 1661 116
rect 1683 119 1685 121
rect 1596 102 1598 104
rect 1740 127 1742 129
rect 1742 119 1744 121
rect 1691 111 1693 113
rect 1772 119 1774 121
rect 1782 132 1784 134
rect 1830 127 1832 129
rect 1813 111 1815 113
rect 1870 136 1872 138
rect 1870 119 1872 121
rect 1902 115 1904 117
rect 1861 111 1863 113
rect 1969 127 1971 129
rect 1925 110 1927 112
rect 2018 127 2020 129
rect 1977 111 1979 113
rect 2058 119 2060 121
rect 2068 132 2070 134
rect 2116 127 2118 129
rect 2099 111 2101 113
rect 2156 136 2158 138
rect 2147 109 2149 111
rect 2156 119 2158 121
rect 2188 115 2190 117
rect 2207 111 2209 113
rect 2236 127 2238 129
rect 2276 111 2278 113
rect 2300 128 2302 130
rect 2276 87 2278 89
rect 2311 83 2313 85
rect 17 59 19 61
rect 41 47 43 49
rect 81 55 83 57
rect 49 39 51 41
rect 89 63 91 65
rect 139 55 141 57
rect 170 55 172 57
rect 133 47 135 49
rect 261 72 263 74
rect 211 63 213 65
rect 180 42 182 44
rect 228 50 230 52
rect 268 61 270 63
rect 268 42 270 44
rect 348 55 350 57
rect 316 39 318 41
rect 291 31 293 33
rect 356 63 358 65
rect 406 55 408 57
rect 437 55 439 57
rect 400 47 402 49
rect 528 72 530 74
rect 478 63 480 65
rect 447 42 449 44
rect 495 50 497 52
rect 535 61 537 63
rect 535 42 537 44
rect 615 55 617 57
rect 583 39 585 41
rect 558 31 560 33
rect 623 63 625 65
rect 673 55 675 57
rect 704 55 706 57
rect 667 47 669 49
rect 795 72 797 74
rect 745 63 747 65
rect 714 42 716 44
rect 762 50 764 52
rect 802 61 804 63
rect 802 42 804 44
rect 882 55 884 57
rect 850 39 852 41
rect 825 31 827 33
rect 890 63 892 65
rect 940 55 942 57
rect 971 55 973 57
rect 934 47 936 49
rect 1062 72 1064 74
rect 1012 63 1014 65
rect 981 42 983 44
rect 1029 50 1031 52
rect 1069 61 1071 63
rect 1069 42 1071 44
rect 1149 55 1151 57
rect 1117 39 1119 41
rect 1092 31 1094 33
rect 1157 63 1159 65
rect 1207 55 1209 57
rect 1238 55 1240 57
rect 1201 47 1203 49
rect 1329 72 1331 74
rect 1279 63 1281 65
rect 1248 42 1250 44
rect 1296 50 1298 52
rect 1336 61 1338 63
rect 1336 42 1338 44
rect 1416 55 1418 57
rect 1384 39 1386 41
rect 1359 31 1361 33
rect 1424 63 1426 65
rect 1474 55 1476 57
rect 1505 55 1507 57
rect 1468 47 1470 49
rect 1596 72 1598 74
rect 1546 63 1548 65
rect 1515 42 1517 44
rect 1563 50 1565 52
rect 1603 61 1605 63
rect 1603 42 1605 44
rect 1683 55 1685 57
rect 1651 39 1653 41
rect 1626 31 1628 33
rect 1691 63 1693 65
rect 1741 55 1743 57
rect 1772 55 1774 57
rect 1735 47 1737 49
rect 1863 72 1865 74
rect 1813 63 1815 65
rect 1782 42 1784 44
rect 1830 50 1832 52
rect 1870 61 1872 63
rect 1870 42 1872 44
rect 1925 64 1927 66
rect 1893 31 1895 33
rect 1969 47 1971 49
rect 1977 63 1979 65
rect 2058 55 2060 57
rect 2018 47 2020 49
rect 2149 72 2151 74
rect 2099 63 2101 65
rect 2068 42 2070 44
rect 2116 50 2118 52
rect 2156 61 2158 63
rect 2156 42 2158 44
rect 2210 63 2212 65
rect 2236 48 2238 50
rect 2180 31 2182 33
rect 2276 63 2278 65
rect 2300 48 2302 50
rect 2320 21 2322 23
rect 9 -14 11 -12
rect 41 -20 43 -18
rect 57 -31 59 -29
rect 81 -25 83 -23
rect 121 -17 123 -15
rect 139 -25 141 -23
rect 89 -33 91 -31
rect 170 -25 172 -23
rect 180 -12 182 -10
rect 227 -17 229 -15
rect 211 -33 213 -31
rect 268 -8 270 -6
rect 259 -33 261 -31
rect 268 -25 270 -23
rect 300 -29 302 -27
rect 324 -31 326 -29
rect 348 -25 350 -23
rect 388 -17 390 -15
rect 406 -25 408 -23
rect 356 -33 358 -31
rect 437 -25 439 -23
rect 447 -12 449 -10
rect 494 -17 496 -15
rect 478 -33 480 -31
rect 535 -8 537 -6
rect 526 -33 528 -31
rect 535 -25 537 -23
rect 567 -29 569 -27
rect 591 -31 593 -29
rect 615 -25 617 -23
rect 655 -17 657 -15
rect 673 -25 675 -23
rect 623 -33 625 -31
rect 704 -25 706 -23
rect 714 -12 716 -10
rect 761 -17 763 -15
rect 745 -33 747 -31
rect 802 -8 804 -6
rect 793 -33 795 -31
rect 802 -25 804 -23
rect 834 -29 836 -27
rect 858 -31 860 -29
rect 882 -25 884 -23
rect 922 -17 924 -15
rect 940 -25 942 -23
rect 890 -33 892 -31
rect 971 -25 973 -23
rect 981 -12 983 -10
rect 1028 -17 1030 -15
rect 1012 -33 1014 -31
rect 1069 -8 1071 -6
rect 1060 -33 1062 -31
rect 1069 -25 1071 -23
rect 1101 -29 1103 -27
rect 1125 -31 1127 -29
rect 1149 -25 1151 -23
rect 1189 -17 1191 -15
rect 1207 -25 1209 -23
rect 1157 -33 1159 -31
rect 1238 -25 1240 -23
rect 1248 -12 1250 -10
rect 1295 -17 1297 -15
rect 1279 -33 1281 -31
rect 1336 -8 1338 -6
rect 1327 -33 1329 -31
rect 1336 -25 1338 -23
rect 1368 -29 1370 -27
rect 1392 -31 1394 -29
rect 1416 -25 1418 -23
rect 1456 -17 1458 -15
rect 1474 -25 1476 -23
rect 1424 -33 1426 -31
rect 1505 -25 1507 -23
rect 1515 -12 1517 -10
rect 1562 -17 1564 -15
rect 1546 -33 1548 -31
rect 1603 -8 1605 -6
rect 1594 -33 1596 -31
rect 1603 -25 1605 -23
rect 1635 -29 1637 -27
rect 1659 -31 1661 -29
rect 1683 -25 1685 -23
rect 1723 -17 1725 -15
rect 1741 -25 1743 -23
rect 1691 -33 1693 -31
rect 1772 -25 1774 -23
rect 1782 -12 1784 -10
rect 1829 -17 1831 -15
rect 1813 -33 1815 -31
rect 1870 -8 1872 -6
rect 1861 -34 1863 -32
rect 1870 -25 1872 -23
rect 1902 -29 1904 -27
rect 1969 -17 1971 -15
rect 1925 -34 1927 -32
rect 2018 -17 2020 -15
rect 1977 -33 1979 -31
rect 2058 -25 2060 -23
rect 2068 -12 2070 -10
rect 2116 -17 2118 -15
rect 2099 -33 2101 -31
rect 2156 -8 2158 -6
rect 2147 -33 2149 -31
rect 2156 -25 2158 -23
rect 2188 -29 2190 -27
rect 2210 -33 2212 -31
rect 2236 -16 2238 -14
rect 2276 -33 2278 -31
rect 2300 -16 2302 -14
rect 2276 -57 2278 -55
rect 2311 -61 2313 -59
rect 17 -85 19 -83
rect 41 -97 43 -95
rect 81 -89 83 -87
rect 49 -105 51 -103
rect 89 -81 91 -79
rect 139 -89 141 -87
rect 170 -89 172 -87
rect 134 -97 136 -95
rect 261 -72 263 -70
rect 211 -81 213 -79
rect 180 -102 182 -100
rect 228 -94 230 -92
rect 268 -83 270 -81
rect 268 -102 270 -100
rect 348 -89 350 -87
rect 316 -105 318 -103
rect 292 -113 294 -111
rect 356 -81 358 -79
rect 406 -89 408 -87
rect 437 -89 439 -87
rect 401 -97 403 -95
rect 528 -72 530 -70
rect 478 -81 480 -79
rect 447 -102 449 -100
rect 495 -94 497 -92
rect 535 -83 537 -81
rect 535 -102 537 -100
rect 615 -89 617 -87
rect 583 -105 585 -103
rect 559 -113 561 -111
rect 623 -81 625 -79
rect 673 -89 675 -87
rect 704 -89 706 -87
rect 668 -97 670 -95
rect 795 -72 797 -70
rect 745 -81 747 -79
rect 714 -102 716 -100
rect 762 -94 764 -92
rect 802 -83 804 -81
rect 802 -102 804 -100
rect 882 -89 884 -87
rect 850 -105 852 -103
rect 826 -113 828 -111
rect 890 -81 892 -79
rect 940 -89 942 -87
rect 971 -89 973 -87
rect 935 -97 937 -95
rect 1062 -72 1064 -70
rect 1012 -81 1014 -79
rect 981 -102 983 -100
rect 1029 -94 1031 -92
rect 1069 -83 1071 -81
rect 1069 -102 1071 -100
rect 1149 -89 1151 -87
rect 1117 -105 1119 -103
rect 1093 -113 1095 -111
rect 1157 -81 1159 -79
rect 1207 -89 1209 -87
rect 1238 -89 1240 -87
rect 1202 -97 1204 -95
rect 1329 -72 1331 -70
rect 1279 -81 1281 -79
rect 1248 -102 1250 -100
rect 1296 -94 1298 -92
rect 1336 -83 1338 -81
rect 1336 -102 1338 -100
rect 1416 -89 1418 -87
rect 1384 -105 1386 -103
rect 1360 -113 1362 -111
rect 1424 -81 1426 -79
rect 1474 -89 1476 -87
rect 1505 -89 1507 -87
rect 1469 -97 1471 -95
rect 1596 -72 1598 -70
rect 1546 -81 1548 -79
rect 1515 -102 1517 -100
rect 1563 -94 1565 -92
rect 1603 -83 1605 -81
rect 1603 -102 1605 -100
rect 1683 -89 1685 -87
rect 1651 -105 1653 -103
rect 1627 -113 1629 -111
rect 1691 -81 1693 -79
rect 1741 -89 1743 -87
rect 1772 -89 1774 -87
rect 1736 -97 1738 -95
rect 1863 -72 1865 -70
rect 1813 -81 1815 -79
rect 1782 -102 1784 -100
rect 1830 -94 1832 -92
rect 1870 -83 1872 -81
rect 1870 -102 1872 -100
rect 1925 -80 1927 -78
rect 1894 -113 1896 -111
rect 1969 -97 1971 -95
rect 1977 -81 1979 -79
rect 2058 -89 2060 -87
rect 2018 -97 2020 -95
rect 2149 -72 2151 -70
rect 2099 -81 2101 -79
rect 2068 -102 2070 -100
rect 2116 -94 2118 -92
rect 2156 -83 2158 -81
rect 2156 -102 2158 -100
rect 2210 -81 2212 -79
rect 2236 -96 2238 -94
rect 2180 -113 2182 -111
rect 2276 -81 2278 -79
rect 2300 -96 2302 -94
rect 2320 -123 2322 -121
rect 9 -158 11 -156
rect 41 -161 43 -159
rect 57 -174 59 -172
rect 81 -169 83 -167
rect 138 -161 140 -159
rect 140 -169 142 -167
rect 89 -177 91 -175
rect 170 -169 172 -167
rect 180 -156 182 -154
rect 228 -161 230 -159
rect 211 -177 213 -175
rect 268 -152 270 -150
rect 268 -169 270 -167
rect 300 -173 302 -171
rect 324 -174 326 -172
rect 348 -169 350 -167
rect 261 -186 263 -184
rect 405 -161 407 -159
rect 407 -169 409 -167
rect 356 -177 358 -175
rect 437 -169 439 -167
rect 447 -156 449 -154
rect 495 -161 497 -159
rect 478 -177 480 -175
rect 535 -152 537 -150
rect 535 -169 537 -167
rect 567 -173 569 -171
rect 591 -174 593 -172
rect 615 -169 617 -167
rect 528 -186 530 -184
rect 672 -161 674 -159
rect 674 -169 676 -167
rect 623 -177 625 -175
rect 704 -169 706 -167
rect 714 -156 716 -154
rect 762 -161 764 -159
rect 745 -177 747 -175
rect 802 -152 804 -150
rect 802 -169 804 -167
rect 834 -173 836 -171
rect 858 -174 860 -172
rect 882 -169 884 -167
rect 795 -186 797 -184
rect 939 -161 941 -159
rect 941 -169 943 -167
rect 890 -177 892 -175
rect 971 -169 973 -167
rect 981 -156 983 -154
rect 1029 -161 1031 -159
rect 1012 -177 1014 -175
rect 1069 -152 1071 -150
rect 1069 -169 1071 -167
rect 1101 -173 1103 -171
rect 1125 -174 1127 -172
rect 1149 -169 1151 -167
rect 1062 -186 1064 -184
rect 1206 -161 1208 -159
rect 1208 -169 1210 -167
rect 1157 -177 1159 -175
rect 1238 -169 1240 -167
rect 1248 -156 1250 -154
rect 1296 -161 1298 -159
rect 1279 -177 1281 -175
rect 1336 -152 1338 -150
rect 1336 -169 1338 -167
rect 1368 -173 1370 -171
rect 1392 -174 1394 -172
rect 1416 -169 1418 -167
rect 1329 -186 1331 -184
rect 1473 -161 1475 -159
rect 1475 -169 1477 -167
rect 1424 -177 1426 -175
rect 1505 -169 1507 -167
rect 1515 -156 1517 -154
rect 1563 -161 1565 -159
rect 1546 -177 1548 -175
rect 1603 -152 1605 -150
rect 1603 -169 1605 -167
rect 1635 -173 1637 -171
rect 1659 -174 1661 -172
rect 1683 -169 1685 -167
rect 1596 -186 1598 -184
rect 1740 -161 1742 -159
rect 1742 -169 1744 -167
rect 1691 -177 1693 -175
rect 1772 -169 1774 -167
rect 1782 -156 1784 -154
rect 1830 -161 1832 -159
rect 1813 -177 1815 -175
rect 1870 -152 1872 -150
rect 1870 -169 1872 -167
rect 1902 -173 1904 -171
rect 1861 -178 1863 -176
rect 1969 -161 1971 -159
rect 1925 -178 1927 -176
rect 2018 -161 2020 -159
rect 1977 -177 1979 -175
rect 2058 -169 2060 -167
rect 2068 -156 2070 -154
rect 2116 -161 2118 -159
rect 2099 -177 2101 -175
rect 2156 -152 2158 -150
rect 2156 -169 2158 -167
rect 2188 -173 2190 -171
rect 2147 -181 2149 -179
rect 2210 -177 2212 -175
rect 2236 -160 2238 -158
rect 2276 -177 2278 -175
rect 2300 -160 2302 -158
rect 2324 -195 2326 -193
rect 2276 -201 2278 -199
rect 133 -204 135 -202
rect 400 -204 402 -202
rect 667 -204 669 -202
rect 934 -204 936 -202
rect 1201 -204 1203 -202
rect 1468 -204 1470 -202
rect 1735 -204 1737 -202
rect 9 -245 11 -243
rect 41 -233 43 -231
rect 49 -246 51 -244
rect 81 -233 83 -231
rect 89 -225 91 -223
rect 139 -233 141 -231
rect 170 -233 172 -231
rect 133 -241 135 -239
rect 261 -216 263 -214
rect 211 -225 213 -223
rect 180 -246 182 -244
rect 228 -238 230 -236
rect 268 -227 270 -225
rect 268 -246 270 -244
rect 316 -246 318 -244
rect 348 -233 350 -231
rect 300 -258 302 -256
rect 356 -225 358 -223
rect 406 -233 408 -231
rect 437 -233 439 -231
rect 400 -241 402 -239
rect 528 -216 530 -214
rect 478 -225 480 -223
rect 447 -246 449 -244
rect 495 -238 497 -236
rect 535 -227 537 -225
rect 535 -246 537 -244
rect 583 -246 585 -244
rect 615 -233 617 -231
rect 567 -258 569 -256
rect 623 -225 625 -223
rect 673 -233 675 -231
rect 704 -233 706 -231
rect 667 -241 669 -239
rect 795 -216 797 -214
rect 745 -225 747 -223
rect 714 -246 716 -244
rect 762 -238 764 -236
rect 802 -227 804 -225
rect 802 -246 804 -244
rect 850 -246 852 -244
rect 882 -233 884 -231
rect 834 -258 836 -256
rect 890 -225 892 -223
rect 940 -233 942 -231
rect 971 -233 973 -231
rect 934 -241 936 -239
rect 1062 -216 1064 -214
rect 1012 -225 1014 -223
rect 981 -246 983 -244
rect 1029 -238 1031 -236
rect 1069 -227 1071 -225
rect 1069 -246 1071 -244
rect 1117 -246 1119 -244
rect 1149 -233 1151 -231
rect 1101 -258 1103 -256
rect 1157 -225 1159 -223
rect 1207 -233 1209 -231
rect 1238 -233 1240 -231
rect 1201 -241 1203 -239
rect 1329 -216 1331 -214
rect 1279 -225 1281 -223
rect 1248 -246 1250 -244
rect 1296 -238 1298 -236
rect 1336 -227 1338 -225
rect 1336 -246 1338 -244
rect 1384 -246 1386 -244
rect 1416 -233 1418 -231
rect 1368 -258 1370 -256
rect 1424 -225 1426 -223
rect 1474 -233 1476 -231
rect 1505 -233 1507 -231
rect 1468 -241 1470 -239
rect 1596 -216 1598 -214
rect 1546 -225 1548 -223
rect 1515 -246 1517 -244
rect 1563 -238 1565 -236
rect 1603 -227 1605 -225
rect 1603 -246 1605 -244
rect 1651 -246 1653 -244
rect 1683 -233 1685 -231
rect 1635 -258 1637 -256
rect 1691 -225 1693 -223
rect 1741 -233 1743 -231
rect 1772 -233 1774 -231
rect 1735 -241 1737 -239
rect 1863 -216 1865 -214
rect 1813 -225 1815 -223
rect 1782 -246 1784 -244
rect 1830 -238 1832 -236
rect 1870 -227 1872 -225
rect 1870 -246 1872 -244
rect 1925 -224 1927 -222
rect 1902 -258 1904 -256
rect 1969 -241 1971 -239
rect 1977 -225 1979 -223
rect 2058 -233 2060 -231
rect 2018 -241 2020 -239
rect 2149 -216 2151 -214
rect 2099 -225 2101 -223
rect 2068 -246 2070 -244
rect 2116 -238 2118 -236
rect 2156 -227 2158 -225
rect 2156 -246 2158 -244
rect 2188 -230 2190 -228
rect 2210 -225 2212 -223
rect 2236 -242 2238 -240
rect 2276 -225 2278 -223
rect 2300 -240 2302 -238
rect 2328 -267 2330 -265
<< via2 >>
rect 2324 301 2326 303
rect 1929 288 1931 290
rect 2092 288 2094 290
rect 3 274 5 276
rect 213 271 215 273
rect 263 272 265 274
rect 352 271 354 273
rect 480 271 482 273
rect 530 271 532 273
rect 619 271 621 273
rect 747 271 749 273
rect 886 271 888 273
rect 1014 271 1016 273
rect 1153 271 1155 273
rect 1281 271 1283 273
rect 1420 271 1422 273
rect 1548 271 1550 273
rect 1687 271 1689 273
rect 1815 271 1817 273
rect 1861 271 1863 273
rect 2092 271 2094 273
rect 2193 271 2195 273
rect 2304 272 2306 274
rect 45 257 47 259
rect 304 259 306 261
rect 312 257 314 259
rect 571 259 573 261
rect 579 257 581 259
rect 838 259 840 261
rect 797 255 799 257
rect 846 257 848 259
rect 1105 259 1107 261
rect 1064 255 1066 257
rect 1113 257 1115 259
rect 1372 259 1374 261
rect 1380 257 1382 259
rect 1639 259 1641 261
rect 1647 257 1649 259
rect 1906 259 1908 261
rect 2192 259 2194 261
rect 1929 254 1931 256
rect 1331 246 1333 248
rect 1598 248 1600 250
rect 213 234 215 236
rect 480 234 482 236
rect 747 234 749 236
rect 1014 234 1016 236
rect 1281 234 1283 236
rect 1548 234 1550 236
rect 1815 234 1817 236
rect 2264 224 2266 226
rect 352 216 354 218
rect 619 216 621 218
rect 886 216 888 218
rect 1153 216 1155 218
rect 1420 216 1422 218
rect 1687 216 1689 218
rect 1881 216 1883 218
rect 3 203 5 205
rect 1929 208 1931 210
rect 2315 227 2317 229
rect 2236 198 2238 200
rect 304 194 306 196
rect 571 194 573 196
rect 838 194 840 196
rect 1105 194 1107 196
rect 1372 194 1374 196
rect 1639 194 1641 196
rect 1906 194 1908 196
rect 2192 194 2194 196
rect 336 191 338 193
rect 603 191 605 193
rect 870 191 872 193
rect 1137 191 1139 193
rect 1404 191 1406 193
rect 1671 191 1673 193
rect 2304 192 2306 194
rect 45 183 47 185
rect 312 183 314 185
rect 579 183 581 185
rect 846 183 848 185
rect 1113 183 1115 185
rect 1380 183 1382 185
rect 1647 183 1649 185
rect 3 130 5 132
rect 2324 165 2326 167
rect 352 127 354 129
rect 619 127 621 129
rect 886 127 888 129
rect 1153 127 1155 129
rect 1420 127 1422 129
rect 1687 127 1689 129
rect 2228 127 2230 129
rect 2304 128 2306 130
rect 45 114 47 116
rect 304 115 306 117
rect 312 114 314 116
rect 571 115 573 117
rect 579 114 581 116
rect 838 115 840 117
rect 846 114 848 116
rect 1105 115 1107 117
rect 1113 114 1115 116
rect 1372 115 1374 117
rect 1380 114 1382 116
rect 1639 115 1641 117
rect 1647 114 1649 116
rect 1906 115 1908 117
rect 2192 115 2194 117
rect 1873 111 1875 113
rect 1929 110 1931 112
rect 336 102 338 104
rect 603 102 605 104
rect 870 102 872 104
rect 1137 102 1139 104
rect 1404 102 1406 104
rect 1671 102 1673 104
rect 1865 77 1867 79
rect 352 72 354 74
rect 619 72 621 74
rect 886 72 888 74
rect 1153 72 1155 74
rect 1420 72 1422 74
rect 1687 72 1689 74
rect 3 59 5 61
rect 1929 64 1931 66
rect 2315 83 2317 85
rect 304 50 306 52
rect 571 50 573 52
rect 838 50 840 52
rect 1105 50 1107 52
rect 1372 50 1374 52
rect 1639 50 1641 52
rect 1906 50 1908 52
rect 2192 50 2194 52
rect 336 47 338 49
rect 603 47 605 49
rect 870 47 872 49
rect 1137 47 1139 49
rect 1404 47 1406 49
rect 1671 47 1673 49
rect 2220 48 2222 50
rect 2304 48 2306 50
rect 45 39 47 41
rect 312 39 314 41
rect 579 39 581 41
rect 846 39 848 41
rect 1113 39 1115 41
rect 1380 39 1382 41
rect 1647 39 1649 41
rect 3 -14 5 -12
rect 2324 21 2326 23
rect 352 -17 354 -15
rect 619 -17 621 -15
rect 886 -17 888 -15
rect 1153 -17 1155 -15
rect 1420 -17 1422 -15
rect 1687 -17 1689 -15
rect 2304 -16 2306 -14
rect 2228 -19 2230 -17
rect 45 -31 47 -29
rect 304 -29 306 -27
rect 312 -31 314 -29
rect 571 -29 573 -27
rect 579 -31 581 -29
rect 838 -29 840 -27
rect 846 -31 848 -29
rect 1105 -29 1107 -27
rect 1113 -31 1115 -29
rect 1372 -29 1374 -27
rect 1380 -31 1382 -29
rect 1639 -29 1641 -27
rect 1647 -31 1649 -29
rect 1906 -29 1908 -27
rect 2192 -29 2194 -27
rect 1857 -34 1859 -32
rect 1929 -34 1931 -32
rect 336 -42 338 -40
rect 603 -42 605 -40
rect 870 -42 872 -40
rect 1137 -42 1139 -40
rect 1404 -42 1406 -40
rect 1671 -42 1673 -40
rect 352 -72 354 -70
rect 619 -72 621 -70
rect 886 -72 888 -70
rect 1153 -72 1155 -70
rect 1420 -72 1422 -70
rect 1687 -72 1689 -70
rect 1849 -72 1851 -70
rect 3 -85 5 -83
rect 1929 -80 1931 -78
rect 2315 -61 2317 -59
rect 304 -94 306 -92
rect 571 -94 573 -92
rect 838 -94 840 -92
rect 1105 -94 1107 -92
rect 1372 -94 1374 -92
rect 1639 -94 1641 -92
rect 1906 -94 1908 -92
rect 2192 -94 2194 -92
rect 336 -97 338 -95
rect 603 -97 605 -95
rect 870 -97 872 -95
rect 1137 -97 1139 -95
rect 1404 -97 1406 -95
rect 1671 -97 1673 -95
rect 2304 -96 2306 -94
rect 2236 -101 2238 -99
rect 45 -105 47 -103
rect 312 -105 314 -103
rect 579 -105 581 -103
rect 846 -105 848 -103
rect 1113 -105 1115 -103
rect 1380 -105 1382 -103
rect 1647 -105 1649 -103
rect 3 -158 5 -156
rect 2324 -123 2326 -121
rect 352 -161 354 -159
rect 619 -161 621 -159
rect 886 -161 888 -159
rect 1153 -161 1155 -159
rect 1420 -161 1422 -159
rect 1687 -161 1689 -159
rect 2308 -160 2310 -158
rect 2196 -164 2198 -162
rect 45 -174 47 -172
rect 304 -173 306 -171
rect 312 -174 314 -172
rect 571 -173 573 -171
rect 579 -174 581 -172
rect 838 -173 840 -171
rect 846 -174 848 -172
rect 1105 -173 1107 -171
rect 1113 -174 1115 -172
rect 1372 -173 1374 -171
rect 1380 -174 1382 -172
rect 1639 -173 1641 -171
rect 1647 -174 1649 -172
rect 1906 -173 1908 -171
rect 2192 -173 2194 -171
rect 1841 -178 1843 -176
rect 1929 -178 1931 -176
rect 336 -186 338 -184
rect 603 -186 605 -184
rect 870 -186 872 -184
rect 1137 -186 1139 -184
rect 1404 -186 1406 -184
rect 1671 -186 1673 -184
rect 2328 -195 2330 -193
rect 129 -204 131 -202
rect 352 -216 354 -214
rect 619 -216 621 -214
rect 886 -216 888 -214
rect 1153 -216 1155 -214
rect 1420 -216 1422 -214
rect 1687 -216 1689 -214
rect 1889 -216 1891 -214
rect 1929 -224 1931 -222
rect 37 -233 39 -231
rect 2200 -230 2202 -228
rect 304 -238 306 -236
rect 571 -238 573 -236
rect 838 -238 840 -236
rect 1105 -238 1107 -236
rect 1372 -238 1374 -236
rect 1639 -238 1641 -236
rect 1906 -238 1908 -236
rect 2192 -238 2194 -236
rect 129 -241 131 -239
rect 396 -241 398 -239
rect 663 -241 665 -239
rect 930 -241 932 -239
rect 1197 -241 1199 -239
rect 1464 -241 1466 -239
rect 1731 -241 1733 -239
rect 2244 -242 2246 -240
rect 2320 -240 2322 -238
rect 3 -245 5 -243
rect 45 -246 47 -244
rect 312 -246 314 -244
rect 579 -246 581 -244
rect 846 -246 848 -244
rect 1113 -246 1115 -244
rect 1380 -246 1382 -244
rect 1647 -246 1649 -244
rect 396 -258 398 -256
rect 663 -258 665 -256
rect 930 -258 932 -256
rect 1197 -258 1199 -256
rect 1464 -258 1466 -256
rect 1731 -258 1733 -256
rect 1897 -258 1899 -256
rect 2328 -271 2330 -269
<< via3 >>
rect 263 284 265 286
rect 530 276 532 278
rect 797 268 799 270
rect 1064 260 1066 262
rect 37 -238 39 -236
rect 1331 252 1333 254
rect 1598 244 1600 246
rect 1861 284 1863 286
rect 1760 -238 1762 -236
rect 1841 -255 1843 -253
rect 1849 -263 1851 -261
rect 1865 -239 1867 -237
rect 1873 -247 1875 -245
rect 2264 301 2266 303
rect 2272 301 2274 303
rect 2280 301 2282 303
rect 2288 301 2290 303
rect 2296 301 2298 303
rect 2304 301 2306 303
rect 2328 301 2330 303
rect 2236 202 2238 204
rect 2315 231 2317 233
rect 2228 135 2230 137
rect 2220 65 2222 67
rect 2212 -19 2214 -17
rect 1881 -255 1883 -253
rect 2204 -101 2206 -99
rect 2196 -156 2198 -154
rect 2328 165 2330 167
rect 2315 87 2317 89
rect 2328 21 2330 23
rect 2315 -57 2317 -55
rect 2328 -123 2330 -121
rect 2312 -160 2314 -158
rect 2328 -207 2330 -205
rect 2244 -229 2246 -227
rect 1889 -263 1891 -261
rect 1857 -271 1859 -269
rect 2334 -271 2336 -269
<< via4 >>
rect 2264 301 2266 303
rect 2272 301 2274 303
rect 2280 301 2282 303
rect 1861 284 1863 286
rect 2244 280 2246 282
rect 2334 301 2336 303
rect 2319 231 2321 233
rect 2334 165 2336 167
rect 2319 87 2321 89
rect 2334 21 2336 23
rect 2319 -57 2321 -55
rect 2334 -123 2336 -121
rect 1849 -255 1851 -253
rect 2324 -207 2326 -205
rect 1857 -263 1859 -261
rect 2334 -267 2336 -265
rect 2280 -271 2282 -269
<< via5 >>
rect 2323 230 2327 234
rect 2323 86 2327 90
rect 2323 -58 2327 -54
rect 2323 -202 2327 -198
<< labels >>
rlabel via1 10 -245 10 -245 1 b0
rlabel via1 10 -156 10 -156 1 b0
rlabel via1 18 -84 18 -84 1 b0
rlabel alu1 10 -8 10 -8 1 b0
rlabel via1 18 60 18 60 1 b0
rlabel via1 10 132 10 132 1 b0
rlabel via1 18 204 18 204 1 b0
rlabel alu1 18 258 18 258 1 a1
rlabel alu1 58 204 58 204 1 a1
rlabel alu1 50 276 50 276 1 a0
rlabel via1 58 258 58 258 1 b1
rlabel alu1 42 -233 42 -233 1 p0
rlabel alu1 18 -228 18 -228 1 a0
rlabel alu1 58 -228 58 -228 1 a7
rlabel alu1 18 -173 18 -173 1 a7
rlabel alu1 50 -156 50 -156 1 a6
rlabel alu1 10 -99 10 -99 1 a6
rlabel alu1 58 -84 58 -84 1 a5
rlabel alu1 18 -30 18 -30 1 a5
rlabel alu1 50 -12 50 -12 1 a4
rlabel alu1 10 43 10 43 1 a4
rlabel alu1 58 60 58 60 1 a3
rlabel alu1 18 115 18 115 1 a3
rlabel alu1 50 132 50 132 1 a2
rlabel alu1 10 189 10 189 1 a2
rlabel alu1 260 269 260 269 1 p1
rlabel via1 325 258 325 258 1 b2
rlabel alu1 317 276 317 276 1 a0
rlabel alu1 325 204 325 204 1 a1
rlabel alu1 317 132 317 132 1 a2
rlabel alu1 325 60 325 60 1 a3
rlabel alu1 317 -12 317 -12 1 a4
rlabel alu1 325 -84 325 -84 1 a5
rlabel alu1 317 -156 317 -156 1 a6
rlabel alu1 325 -228 325 -228 1 a7
rlabel alu1 527 269 527 269 1 p2
rlabel alu1 584 276 584 276 1 a0
rlabel alu1 592 204 592 204 1 a1
rlabel alu1 584 132 584 132 1 a2
rlabel alu1 592 60 592 60 1 a3
rlabel alu1 584 -12 584 -12 1 a4
rlabel alu1 592 -84 592 -84 1 a5
rlabel alu1 584 -156 584 -156 1 a6
rlabel alu1 592 -228 592 -228 1 a7
rlabel via1 592 258 592 258 1 b3
rlabel alu1 794 269 794 269 1 p3
rlabel alu1 851 276 851 276 1 a0
rlabel alu1 859 204 859 204 1 a1
rlabel alu1 851 132 851 132 1 a2
rlabel alu1 859 60 859 60 1 a3
rlabel alu1 851 -12 851 -12 1 a4
rlabel alu1 859 -84 859 -84 1 a5
rlabel alu1 851 -156 851 -156 1 a6
rlabel alu1 859 -228 859 -228 1 a7
rlabel via1 859 258 859 258 1 b4
rlabel alu1 1061 269 1061 269 1 p4
rlabel via1 1126 258 1126 258 1 b5
rlabel alu1 1118 276 1118 276 1 a0
rlabel alu1 1118 132 1118 132 1 a2
rlabel alu1 1126 204 1126 204 1 a1
rlabel alu1 1126 60 1126 60 1 a3
rlabel alu1 1118 -12 1118 -12 1 a4
rlabel alu1 1126 -84 1126 -84 1 a5
rlabel alu1 1118 -156 1118 -156 1 a6
rlabel alu1 1126 -228 1126 -228 1 a7
rlabel alu1 1328 269 1328 269 1 p5
rlabel alu1 1385 276 1385 276 1 a0
rlabel via1 1393 258 1393 258 1 b6
rlabel alu1 1393 204 1393 204 1 a1
rlabel alu1 1385 132 1385 132 1 a2
rlabel alu1 1393 60 1393 60 1 a3
rlabel alu1 1385 -12 1385 -12 1 a4
rlabel alu1 1393 -84 1393 -84 1 a5
rlabel alu1 1385 -156 1385 -156 1 a6
rlabel alu1 1393 -228 1393 -228 1 a7
rlabel alu1 1595 269 1595 269 1 p6
rlabel alu1 1652 276 1652 276 1 a0
rlabel via1 1660 258 1660 258 1 b7
rlabel alu1 1660 204 1660 204 1 a1
rlabel alu1 1652 132 1652 132 1 a2
rlabel alu1 1660 60 1660 60 1 a3
rlabel alu1 1652 -12 1652 -12 1 a4
rlabel alu1 1660 -84 1660 -84 1 a5
rlabel alu1 1652 -156 1652 -156 1 a6
rlabel alu1 1660 -228 1660 -228 1 a7
rlabel alu1 1862 -232 1862 -232 1 p14
rlabel alu1 1862 -163 1862 -163 1 p13
rlabel alu1 1862 -88 1862 -88 1 p12
rlabel alu1 1862 -19 1862 -19 1 p11
rlabel alu1 1862 56 1862 56 1 p10
rlabel alu1 1862 125 1862 125 1 p9
rlabel alu1 1862 200 1862 200 1 p8
rlabel alu1 1862 269 1862 269 1 p7
rlabel alu1 1903 -229 1903 -229 1 p15
rlabel alu1 2148 -231 2148 -231 1 s7
rlabel alu1 2148 -173 2148 -173 1 s6
rlabel alu1 2148 -86 2148 -86 1 s5
rlabel alu1 2148 -28 2148 -28 1 s4
rlabel alu1 2148 58 2148 58 1 s3
rlabel alu1 2148 113 2148 113 1 s2
rlabel alu1 2148 201 2148 201 1 s1
rlabel alu1 2148 269 2148 269 1 s0
rlabel alu1 1915 287 1915 287 1 b0
rlabel alu1 1915 176 1915 176 1 b1
rlabel alu1 1915 144 1915 144 1 b2
rlabel alu1 1915 32 1915 32 1 b3
rlabel alu1 1915 -1 1915 -1 1 b4
rlabel alu1 1915 -112 1915 -112 1 b5
rlabel alu1 1915 -144 1915 -144 1 b6
rlabel alu1 1915 -255 1915 -255 1 b7
rlabel alu1 2034 264 2034 264 1 a0
rlabel alu1 2034 200 2034 200 1 a1
rlabel alu1 2034 120 2034 120 1 a2
rlabel alu1 2034 56 2034 56 1 a3
rlabel alu1 2034 -24 2034 -24 1 a4
rlabel alu1 2034 -88 2034 -88 1 a5
rlabel alu1 2034 -168 2034 -168 1 a6
rlabel alu1 2034 -232 2034 -232 1 a7
rlabel alu1 2257 264 2257 264 1 out0
rlabel alu1 2257 200 2257 200 1 out1
rlabel alu1 2257 120 2257 120 1 out2
rlabel alu1 2257 56 2257 56 1 out3
rlabel alu1 2257 -24 2257 -24 1 out4
rlabel alu1 2257 -88 2257 -88 1 out5
rlabel alu1 2257 -168 2257 -168 1 out6
rlabel alu1 2257 -232 2257 -232 1 out7
rlabel alu1 2325 264 2325 264 1 out8
rlabel alu1 2325 200 2325 200 1 out9
rlabel alu1 2325 120 2325 120 1 out10
rlabel alu1 2325 56 2325 56 1 out11
rlabel alu1 2325 -24 2325 -24 1 out12
rlabel alu1 2325 -88 2325 -88 1 out13
rlabel alu1 2325 -168 2325 -168 1 out14
rlabel alu1 2325 -232 2325 -232 1 out15
rlabel alu5 2337 314 2337 314 1 Vdd
rlabel alu6 2346 314 2346 314 7 Gnd
rlabel alu1 1923 256 1923 256 1 cin
rlabel alu1 1923 208 1923 208 1 cin
rlabel alu1 1923 112 1923 112 1 cin
rlabel alu1 1923 64 1923 64 1 cin
rlabel alu1 1923 -32 1923 -32 1 cin
rlabel alu1 1923 -80 1923 -80 1 cin
rlabel alu2 1924 -176 1924 -176 1 cin
rlabel alu2 1924 -224 1924 -224 1 cin
rlabel alu1 2201 -258 2201 -258 1 sel
rlabel alu1 2269 -258 2269 -258 1 sel
rlabel alu1 2201 -144 2201 -144 1 sel
rlabel alu1 2269 -144 2269 -144 1 sel
rlabel alu1 2201 -112 2201 -112 1 sel
rlabel alu1 2269 -112 2269 -112 1 sel
rlabel alu1 2201 0 2201 0 1 sel
rlabel alu1 2269 0 2269 0 1 sel
rlabel alu1 2201 32 2201 32 1 sel
rlabel alu1 2269 32 2269 32 1 sel
rlabel alu1 2201 144 2201 144 1 sel
rlabel alu1 2269 144 2269 144 1 sel
rlabel alu1 2201 176 2201 176 1 sel
rlabel alu1 2269 176 2269 176 1 sel
rlabel alu1 2201 288 2201 288 1 sel
rlabel alu1 2269 288 2269 288 1 sel
<< end >>
